magic
tech sky130A
magscale 1 2
timestamp 1713233265
<< pwell >>
rect -2521 -1058 2521 1058
<< mvnmos >>
rect -2293 -800 -2093 800
rect -2035 -800 -1835 800
rect -1777 -800 -1577 800
rect -1519 -800 -1319 800
rect -1261 -800 -1061 800
rect -1003 -800 -803 800
rect -745 -800 -545 800
rect -487 -800 -287 800
rect -229 -800 -29 800
rect 29 -800 229 800
rect 287 -800 487 800
rect 545 -800 745 800
rect 803 -800 1003 800
rect 1061 -800 1261 800
rect 1319 -800 1519 800
rect 1577 -800 1777 800
rect 1835 -800 2035 800
rect 2093 -800 2293 800
<< mvndiff >>
rect -2351 788 -2293 800
rect -2351 -788 -2339 788
rect -2305 -788 -2293 788
rect -2351 -800 -2293 -788
rect -2093 788 -2035 800
rect -2093 -788 -2081 788
rect -2047 -788 -2035 788
rect -2093 -800 -2035 -788
rect -1835 788 -1777 800
rect -1835 -788 -1823 788
rect -1789 -788 -1777 788
rect -1835 -800 -1777 -788
rect -1577 788 -1519 800
rect -1577 -788 -1565 788
rect -1531 -788 -1519 788
rect -1577 -800 -1519 -788
rect -1319 788 -1261 800
rect -1319 -788 -1307 788
rect -1273 -788 -1261 788
rect -1319 -800 -1261 -788
rect -1061 788 -1003 800
rect -1061 -788 -1049 788
rect -1015 -788 -1003 788
rect -1061 -800 -1003 -788
rect -803 788 -745 800
rect -803 -788 -791 788
rect -757 -788 -745 788
rect -803 -800 -745 -788
rect -545 788 -487 800
rect -545 -788 -533 788
rect -499 -788 -487 788
rect -545 -800 -487 -788
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
rect 487 788 545 800
rect 487 -788 499 788
rect 533 -788 545 788
rect 487 -800 545 -788
rect 745 788 803 800
rect 745 -788 757 788
rect 791 -788 803 788
rect 745 -800 803 -788
rect 1003 788 1061 800
rect 1003 -788 1015 788
rect 1049 -788 1061 788
rect 1003 -800 1061 -788
rect 1261 788 1319 800
rect 1261 -788 1273 788
rect 1307 -788 1319 788
rect 1261 -800 1319 -788
rect 1519 788 1577 800
rect 1519 -788 1531 788
rect 1565 -788 1577 788
rect 1519 -800 1577 -788
rect 1777 788 1835 800
rect 1777 -788 1789 788
rect 1823 -788 1835 788
rect 1777 -800 1835 -788
rect 2035 788 2093 800
rect 2035 -788 2047 788
rect 2081 -788 2093 788
rect 2035 -800 2093 -788
rect 2293 788 2351 800
rect 2293 -788 2305 788
rect 2339 -788 2351 788
rect 2293 -800 2351 -788
<< mvndiffc >>
rect -2339 -788 -2305 788
rect -2081 -788 -2047 788
rect -1823 -788 -1789 788
rect -1565 -788 -1531 788
rect -1307 -788 -1273 788
rect -1049 -788 -1015 788
rect -791 -788 -757 788
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
rect 757 -788 791 788
rect 1015 -788 1049 788
rect 1273 -788 1307 788
rect 1531 -788 1565 788
rect 1789 -788 1823 788
rect 2047 -788 2081 788
rect 2305 -788 2339 788
<< mvpsubdiff >>
rect -2485 1010 2485 1022
rect -2485 976 -2377 1010
rect 2377 976 2485 1010
rect -2485 964 2485 976
rect -2485 914 -2427 964
rect -2485 -914 -2473 914
rect -2439 -914 -2427 914
rect 2427 914 2485 964
rect -2485 -964 -2427 -914
rect 2427 -914 2439 914
rect 2473 -914 2485 914
rect 2427 -964 2485 -914
rect -2485 -976 2485 -964
rect -2485 -1010 -2377 -976
rect 2377 -1010 2485 -976
rect -2485 -1022 2485 -1010
<< mvpsubdiffcont >>
rect -2377 976 2377 1010
rect -2473 -914 -2439 914
rect 2439 -914 2473 914
rect -2377 -1010 2377 -976
<< poly >>
rect -2293 872 -2093 888
rect -2293 838 -2277 872
rect -2109 838 -2093 872
rect -2293 800 -2093 838
rect -2035 872 -1835 888
rect -2035 838 -2019 872
rect -1851 838 -1835 872
rect -2035 800 -1835 838
rect -1777 872 -1577 888
rect -1777 838 -1761 872
rect -1593 838 -1577 872
rect -1777 800 -1577 838
rect -1519 872 -1319 888
rect -1519 838 -1503 872
rect -1335 838 -1319 872
rect -1519 800 -1319 838
rect -1261 872 -1061 888
rect -1261 838 -1245 872
rect -1077 838 -1061 872
rect -1261 800 -1061 838
rect -1003 872 -803 888
rect -1003 838 -987 872
rect -819 838 -803 872
rect -1003 800 -803 838
rect -745 872 -545 888
rect -745 838 -729 872
rect -561 838 -545 872
rect -745 800 -545 838
rect -487 872 -287 888
rect -487 838 -471 872
rect -303 838 -287 872
rect -487 800 -287 838
rect -229 872 -29 888
rect -229 838 -213 872
rect -45 838 -29 872
rect -229 800 -29 838
rect 29 872 229 888
rect 29 838 45 872
rect 213 838 229 872
rect 29 800 229 838
rect 287 872 487 888
rect 287 838 303 872
rect 471 838 487 872
rect 287 800 487 838
rect 545 872 745 888
rect 545 838 561 872
rect 729 838 745 872
rect 545 800 745 838
rect 803 872 1003 888
rect 803 838 819 872
rect 987 838 1003 872
rect 803 800 1003 838
rect 1061 872 1261 888
rect 1061 838 1077 872
rect 1245 838 1261 872
rect 1061 800 1261 838
rect 1319 872 1519 888
rect 1319 838 1335 872
rect 1503 838 1519 872
rect 1319 800 1519 838
rect 1577 872 1777 888
rect 1577 838 1593 872
rect 1761 838 1777 872
rect 1577 800 1777 838
rect 1835 872 2035 888
rect 1835 838 1851 872
rect 2019 838 2035 872
rect 1835 800 2035 838
rect 2093 872 2293 888
rect 2093 838 2109 872
rect 2277 838 2293 872
rect 2093 800 2293 838
rect -2293 -838 -2093 -800
rect -2293 -872 -2277 -838
rect -2109 -872 -2093 -838
rect -2293 -888 -2093 -872
rect -2035 -838 -1835 -800
rect -2035 -872 -2019 -838
rect -1851 -872 -1835 -838
rect -2035 -888 -1835 -872
rect -1777 -838 -1577 -800
rect -1777 -872 -1761 -838
rect -1593 -872 -1577 -838
rect -1777 -888 -1577 -872
rect -1519 -838 -1319 -800
rect -1519 -872 -1503 -838
rect -1335 -872 -1319 -838
rect -1519 -888 -1319 -872
rect -1261 -838 -1061 -800
rect -1261 -872 -1245 -838
rect -1077 -872 -1061 -838
rect -1261 -888 -1061 -872
rect -1003 -838 -803 -800
rect -1003 -872 -987 -838
rect -819 -872 -803 -838
rect -1003 -888 -803 -872
rect -745 -838 -545 -800
rect -745 -872 -729 -838
rect -561 -872 -545 -838
rect -745 -888 -545 -872
rect -487 -838 -287 -800
rect -487 -872 -471 -838
rect -303 -872 -287 -838
rect -487 -888 -287 -872
rect -229 -838 -29 -800
rect -229 -872 -213 -838
rect -45 -872 -29 -838
rect -229 -888 -29 -872
rect 29 -838 229 -800
rect 29 -872 45 -838
rect 213 -872 229 -838
rect 29 -888 229 -872
rect 287 -838 487 -800
rect 287 -872 303 -838
rect 471 -872 487 -838
rect 287 -888 487 -872
rect 545 -838 745 -800
rect 545 -872 561 -838
rect 729 -872 745 -838
rect 545 -888 745 -872
rect 803 -838 1003 -800
rect 803 -872 819 -838
rect 987 -872 1003 -838
rect 803 -888 1003 -872
rect 1061 -838 1261 -800
rect 1061 -872 1077 -838
rect 1245 -872 1261 -838
rect 1061 -888 1261 -872
rect 1319 -838 1519 -800
rect 1319 -872 1335 -838
rect 1503 -872 1519 -838
rect 1319 -888 1519 -872
rect 1577 -838 1777 -800
rect 1577 -872 1593 -838
rect 1761 -872 1777 -838
rect 1577 -888 1777 -872
rect 1835 -838 2035 -800
rect 1835 -872 1851 -838
rect 2019 -872 2035 -838
rect 1835 -888 2035 -872
rect 2093 -838 2293 -800
rect 2093 -872 2109 -838
rect 2277 -872 2293 -838
rect 2093 -888 2293 -872
<< polycont >>
rect -2277 838 -2109 872
rect -2019 838 -1851 872
rect -1761 838 -1593 872
rect -1503 838 -1335 872
rect -1245 838 -1077 872
rect -987 838 -819 872
rect -729 838 -561 872
rect -471 838 -303 872
rect -213 838 -45 872
rect 45 838 213 872
rect 303 838 471 872
rect 561 838 729 872
rect 819 838 987 872
rect 1077 838 1245 872
rect 1335 838 1503 872
rect 1593 838 1761 872
rect 1851 838 2019 872
rect 2109 838 2277 872
rect -2277 -872 -2109 -838
rect -2019 -872 -1851 -838
rect -1761 -872 -1593 -838
rect -1503 -872 -1335 -838
rect -1245 -872 -1077 -838
rect -987 -872 -819 -838
rect -729 -872 -561 -838
rect -471 -872 -303 -838
rect -213 -872 -45 -838
rect 45 -872 213 -838
rect 303 -872 471 -838
rect 561 -872 729 -838
rect 819 -872 987 -838
rect 1077 -872 1245 -838
rect 1335 -872 1503 -838
rect 1593 -872 1761 -838
rect 1851 -872 2019 -838
rect 2109 -872 2277 -838
<< locali >>
rect -2473 976 -2377 1010
rect 2377 976 2473 1010
rect -2473 914 -2439 976
rect 2439 914 2473 976
rect -2293 838 -2277 872
rect -2109 838 -2093 872
rect -2035 838 -2019 872
rect -1851 838 -1835 872
rect -1777 838 -1761 872
rect -1593 838 -1577 872
rect -1519 838 -1503 872
rect -1335 838 -1319 872
rect -1261 838 -1245 872
rect -1077 838 -1061 872
rect -1003 838 -987 872
rect -819 838 -803 872
rect -745 838 -729 872
rect -561 838 -545 872
rect -487 838 -471 872
rect -303 838 -287 872
rect -229 838 -213 872
rect -45 838 -29 872
rect 29 838 45 872
rect 213 838 229 872
rect 287 838 303 872
rect 471 838 487 872
rect 545 838 561 872
rect 729 838 745 872
rect 803 838 819 872
rect 987 838 1003 872
rect 1061 838 1077 872
rect 1245 838 1261 872
rect 1319 838 1335 872
rect 1503 838 1519 872
rect 1577 838 1593 872
rect 1761 838 1777 872
rect 1835 838 1851 872
rect 2019 838 2035 872
rect 2093 838 2109 872
rect 2277 838 2293 872
rect -2339 788 -2305 804
rect -2339 -804 -2305 -788
rect -2081 788 -2047 804
rect -2081 -804 -2047 -788
rect -1823 788 -1789 804
rect -1823 -804 -1789 -788
rect -1565 788 -1531 804
rect -1565 -804 -1531 -788
rect -1307 788 -1273 804
rect -1307 -804 -1273 -788
rect -1049 788 -1015 804
rect -1049 -804 -1015 -788
rect -791 788 -757 804
rect -791 -804 -757 -788
rect -533 788 -499 804
rect -533 -804 -499 -788
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
rect 499 788 533 804
rect 499 -804 533 -788
rect 757 788 791 804
rect 757 -804 791 -788
rect 1015 788 1049 804
rect 1015 -804 1049 -788
rect 1273 788 1307 804
rect 1273 -804 1307 -788
rect 1531 788 1565 804
rect 1531 -804 1565 -788
rect 1789 788 1823 804
rect 1789 -804 1823 -788
rect 2047 788 2081 804
rect 2047 -804 2081 -788
rect 2305 788 2339 804
rect 2305 -804 2339 -788
rect -2293 -872 -2277 -838
rect -2109 -872 -2093 -838
rect -2035 -872 -2019 -838
rect -1851 -872 -1835 -838
rect -1777 -872 -1761 -838
rect -1593 -872 -1577 -838
rect -1519 -872 -1503 -838
rect -1335 -872 -1319 -838
rect -1261 -872 -1245 -838
rect -1077 -872 -1061 -838
rect -1003 -872 -987 -838
rect -819 -872 -803 -838
rect -745 -872 -729 -838
rect -561 -872 -545 -838
rect -487 -872 -471 -838
rect -303 -872 -287 -838
rect -229 -872 -213 -838
rect -45 -872 -29 -838
rect 29 -872 45 -838
rect 213 -872 229 -838
rect 287 -872 303 -838
rect 471 -872 487 -838
rect 545 -872 561 -838
rect 729 -872 745 -838
rect 803 -872 819 -838
rect 987 -872 1003 -838
rect 1061 -872 1077 -838
rect 1245 -872 1261 -838
rect 1319 -872 1335 -838
rect 1503 -872 1519 -838
rect 1577 -872 1593 -838
rect 1761 -872 1777 -838
rect 1835 -872 1851 -838
rect 2019 -872 2035 -838
rect 2093 -872 2109 -838
rect 2277 -872 2293 -838
rect -2473 -976 -2439 -914
rect 2439 -976 2473 -914
rect -2473 -1010 -2377 -976
rect 2377 -1010 2473 -976
<< viali >>
rect -2277 838 -2109 872
rect -2019 838 -1851 872
rect -1761 838 -1593 872
rect -1503 838 -1335 872
rect -1245 838 -1077 872
rect -987 838 -819 872
rect -729 838 -561 872
rect -471 838 -303 872
rect -213 838 -45 872
rect 45 838 213 872
rect 303 838 471 872
rect 561 838 729 872
rect 819 838 987 872
rect 1077 838 1245 872
rect 1335 838 1503 872
rect 1593 838 1761 872
rect 1851 838 2019 872
rect 2109 838 2277 872
rect -2339 -788 -2305 788
rect -2081 -788 -2047 788
rect -1823 -788 -1789 788
rect -1565 -788 -1531 788
rect -1307 -788 -1273 788
rect -1049 -788 -1015 788
rect -791 -788 -757 788
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
rect 757 -788 791 788
rect 1015 -788 1049 788
rect 1273 -788 1307 788
rect 1531 -788 1565 788
rect 1789 -788 1823 788
rect 2047 -788 2081 788
rect 2305 -788 2339 788
rect -2277 -872 -2109 -838
rect -2019 -872 -1851 -838
rect -1761 -872 -1593 -838
rect -1503 -872 -1335 -838
rect -1245 -872 -1077 -838
rect -987 -872 -819 -838
rect -729 -872 -561 -838
rect -471 -872 -303 -838
rect -213 -872 -45 -838
rect 45 -872 213 -838
rect 303 -872 471 -838
rect 561 -872 729 -838
rect 819 -872 987 -838
rect 1077 -872 1245 -838
rect 1335 -872 1503 -838
rect 1593 -872 1761 -838
rect 1851 -872 2019 -838
rect 2109 -872 2277 -838
<< metal1 >>
rect -2289 872 -2097 878
rect -2289 838 -2277 872
rect -2109 838 -2097 872
rect -2289 832 -2097 838
rect -2031 872 -1839 878
rect -2031 838 -2019 872
rect -1851 838 -1839 872
rect -2031 832 -1839 838
rect -1773 872 -1581 878
rect -1773 838 -1761 872
rect -1593 838 -1581 872
rect -1773 832 -1581 838
rect -1515 872 -1323 878
rect -1515 838 -1503 872
rect -1335 838 -1323 872
rect -1515 832 -1323 838
rect -1257 872 -1065 878
rect -1257 838 -1245 872
rect -1077 838 -1065 872
rect -1257 832 -1065 838
rect -999 872 -807 878
rect -999 838 -987 872
rect -819 838 -807 872
rect -999 832 -807 838
rect -741 872 -549 878
rect -741 838 -729 872
rect -561 838 -549 872
rect -741 832 -549 838
rect -483 872 -291 878
rect -483 838 -471 872
rect -303 838 -291 872
rect -483 832 -291 838
rect -225 872 -33 878
rect -225 838 -213 872
rect -45 838 -33 872
rect -225 832 -33 838
rect 33 872 225 878
rect 33 838 45 872
rect 213 838 225 872
rect 33 832 225 838
rect 291 872 483 878
rect 291 838 303 872
rect 471 838 483 872
rect 291 832 483 838
rect 549 872 741 878
rect 549 838 561 872
rect 729 838 741 872
rect 549 832 741 838
rect 807 872 999 878
rect 807 838 819 872
rect 987 838 999 872
rect 807 832 999 838
rect 1065 872 1257 878
rect 1065 838 1077 872
rect 1245 838 1257 872
rect 1065 832 1257 838
rect 1323 872 1515 878
rect 1323 838 1335 872
rect 1503 838 1515 872
rect 1323 832 1515 838
rect 1581 872 1773 878
rect 1581 838 1593 872
rect 1761 838 1773 872
rect 1581 832 1773 838
rect 1839 872 2031 878
rect 1839 838 1851 872
rect 2019 838 2031 872
rect 1839 832 2031 838
rect 2097 872 2289 878
rect 2097 838 2109 872
rect 2277 838 2289 872
rect 2097 832 2289 838
rect -2345 788 -2299 800
rect -2345 -788 -2339 788
rect -2305 -788 -2299 788
rect -2345 -800 -2299 -788
rect -2087 788 -2041 800
rect -2087 -788 -2081 788
rect -2047 -788 -2041 788
rect -2087 -800 -2041 -788
rect -1829 788 -1783 800
rect -1829 -788 -1823 788
rect -1789 -788 -1783 788
rect -1829 -800 -1783 -788
rect -1571 788 -1525 800
rect -1571 -788 -1565 788
rect -1531 -788 -1525 788
rect -1571 -800 -1525 -788
rect -1313 788 -1267 800
rect -1313 -788 -1307 788
rect -1273 -788 -1267 788
rect -1313 -800 -1267 -788
rect -1055 788 -1009 800
rect -1055 -788 -1049 788
rect -1015 -788 -1009 788
rect -1055 -800 -1009 -788
rect -797 788 -751 800
rect -797 -788 -791 788
rect -757 -788 -751 788
rect -797 -800 -751 -788
rect -539 788 -493 800
rect -539 -788 -533 788
rect -499 -788 -493 788
rect -539 -800 -493 -788
rect -281 788 -235 800
rect -281 -788 -275 788
rect -241 -788 -235 788
rect -281 -800 -235 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 235 788 281 800
rect 235 -788 241 788
rect 275 -788 281 788
rect 235 -800 281 -788
rect 493 788 539 800
rect 493 -788 499 788
rect 533 -788 539 788
rect 493 -800 539 -788
rect 751 788 797 800
rect 751 -788 757 788
rect 791 -788 797 788
rect 751 -800 797 -788
rect 1009 788 1055 800
rect 1009 -788 1015 788
rect 1049 -788 1055 788
rect 1009 -800 1055 -788
rect 1267 788 1313 800
rect 1267 -788 1273 788
rect 1307 -788 1313 788
rect 1267 -800 1313 -788
rect 1525 788 1571 800
rect 1525 -788 1531 788
rect 1565 -788 1571 788
rect 1525 -800 1571 -788
rect 1783 788 1829 800
rect 1783 -788 1789 788
rect 1823 -788 1829 788
rect 1783 -800 1829 -788
rect 2041 788 2087 800
rect 2041 -788 2047 788
rect 2081 -788 2087 788
rect 2041 -800 2087 -788
rect 2299 788 2345 800
rect 2299 -788 2305 788
rect 2339 -788 2345 788
rect 2299 -800 2345 -788
rect -2289 -838 -2097 -832
rect -2289 -872 -2277 -838
rect -2109 -872 -2097 -838
rect -2289 -878 -2097 -872
rect -2031 -838 -1839 -832
rect -2031 -872 -2019 -838
rect -1851 -872 -1839 -838
rect -2031 -878 -1839 -872
rect -1773 -838 -1581 -832
rect -1773 -872 -1761 -838
rect -1593 -872 -1581 -838
rect -1773 -878 -1581 -872
rect -1515 -838 -1323 -832
rect -1515 -872 -1503 -838
rect -1335 -872 -1323 -838
rect -1515 -878 -1323 -872
rect -1257 -838 -1065 -832
rect -1257 -872 -1245 -838
rect -1077 -872 -1065 -838
rect -1257 -878 -1065 -872
rect -999 -838 -807 -832
rect -999 -872 -987 -838
rect -819 -872 -807 -838
rect -999 -878 -807 -872
rect -741 -838 -549 -832
rect -741 -872 -729 -838
rect -561 -872 -549 -838
rect -741 -878 -549 -872
rect -483 -838 -291 -832
rect -483 -872 -471 -838
rect -303 -872 -291 -838
rect -483 -878 -291 -872
rect -225 -838 -33 -832
rect -225 -872 -213 -838
rect -45 -872 -33 -838
rect -225 -878 -33 -872
rect 33 -838 225 -832
rect 33 -872 45 -838
rect 213 -872 225 -838
rect 33 -878 225 -872
rect 291 -838 483 -832
rect 291 -872 303 -838
rect 471 -872 483 -838
rect 291 -878 483 -872
rect 549 -838 741 -832
rect 549 -872 561 -838
rect 729 -872 741 -838
rect 549 -878 741 -872
rect 807 -838 999 -832
rect 807 -872 819 -838
rect 987 -872 999 -838
rect 807 -878 999 -872
rect 1065 -838 1257 -832
rect 1065 -872 1077 -838
rect 1245 -872 1257 -838
rect 1065 -878 1257 -872
rect 1323 -838 1515 -832
rect 1323 -872 1335 -838
rect 1503 -872 1515 -838
rect 1323 -878 1515 -872
rect 1581 -838 1773 -832
rect 1581 -872 1593 -838
rect 1761 -872 1773 -838
rect 1581 -878 1773 -872
rect 1839 -838 2031 -832
rect 1839 -872 1851 -838
rect 2019 -872 2031 -838
rect 1839 -878 2031 -872
rect 2097 -838 2289 -832
rect 2097 -872 2109 -838
rect 2277 -872 2289 -838
rect 2097 -878 2289 -872
<< properties >>
string FIXED_BBOX -2456 -993 2456 993
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 1 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

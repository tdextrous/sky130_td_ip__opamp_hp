magic
tech sky130A
magscale 1 2
timestamp 1713234499
<< nwell >>
rect -2551 -1897 2551 1897
<< mvpmos >>
rect -2293 -1600 -2093 1600
rect -2035 -1600 -1835 1600
rect -1777 -1600 -1577 1600
rect -1519 -1600 -1319 1600
rect -1261 -1600 -1061 1600
rect -1003 -1600 -803 1600
rect -745 -1600 -545 1600
rect -487 -1600 -287 1600
rect -229 -1600 -29 1600
rect 29 -1600 229 1600
rect 287 -1600 487 1600
rect 545 -1600 745 1600
rect 803 -1600 1003 1600
rect 1061 -1600 1261 1600
rect 1319 -1600 1519 1600
rect 1577 -1600 1777 1600
rect 1835 -1600 2035 1600
rect 2093 -1600 2293 1600
<< mvpdiff >>
rect -2351 1588 -2293 1600
rect -2351 -1588 -2339 1588
rect -2305 -1588 -2293 1588
rect -2351 -1600 -2293 -1588
rect -2093 1588 -2035 1600
rect -2093 -1588 -2081 1588
rect -2047 -1588 -2035 1588
rect -2093 -1600 -2035 -1588
rect -1835 1588 -1777 1600
rect -1835 -1588 -1823 1588
rect -1789 -1588 -1777 1588
rect -1835 -1600 -1777 -1588
rect -1577 1588 -1519 1600
rect -1577 -1588 -1565 1588
rect -1531 -1588 -1519 1588
rect -1577 -1600 -1519 -1588
rect -1319 1588 -1261 1600
rect -1319 -1588 -1307 1588
rect -1273 -1588 -1261 1588
rect -1319 -1600 -1261 -1588
rect -1061 1588 -1003 1600
rect -1061 -1588 -1049 1588
rect -1015 -1588 -1003 1588
rect -1061 -1600 -1003 -1588
rect -803 1588 -745 1600
rect -803 -1588 -791 1588
rect -757 -1588 -745 1588
rect -803 -1600 -745 -1588
rect -545 1588 -487 1600
rect -545 -1588 -533 1588
rect -499 -1588 -487 1588
rect -545 -1600 -487 -1588
rect -287 1588 -229 1600
rect -287 -1588 -275 1588
rect -241 -1588 -229 1588
rect -287 -1600 -229 -1588
rect -29 1588 29 1600
rect -29 -1588 -17 1588
rect 17 -1588 29 1588
rect -29 -1600 29 -1588
rect 229 1588 287 1600
rect 229 -1588 241 1588
rect 275 -1588 287 1588
rect 229 -1600 287 -1588
rect 487 1588 545 1600
rect 487 -1588 499 1588
rect 533 -1588 545 1588
rect 487 -1600 545 -1588
rect 745 1588 803 1600
rect 745 -1588 757 1588
rect 791 -1588 803 1588
rect 745 -1600 803 -1588
rect 1003 1588 1061 1600
rect 1003 -1588 1015 1588
rect 1049 -1588 1061 1588
rect 1003 -1600 1061 -1588
rect 1261 1588 1319 1600
rect 1261 -1588 1273 1588
rect 1307 -1588 1319 1588
rect 1261 -1600 1319 -1588
rect 1519 1588 1577 1600
rect 1519 -1588 1531 1588
rect 1565 -1588 1577 1588
rect 1519 -1600 1577 -1588
rect 1777 1588 1835 1600
rect 1777 -1588 1789 1588
rect 1823 -1588 1835 1588
rect 1777 -1600 1835 -1588
rect 2035 1588 2093 1600
rect 2035 -1588 2047 1588
rect 2081 -1588 2093 1588
rect 2035 -1600 2093 -1588
rect 2293 1588 2351 1600
rect 2293 -1588 2305 1588
rect 2339 -1588 2351 1588
rect 2293 -1600 2351 -1588
<< mvpdiffc >>
rect -2339 -1588 -2305 1588
rect -2081 -1588 -2047 1588
rect -1823 -1588 -1789 1588
rect -1565 -1588 -1531 1588
rect -1307 -1588 -1273 1588
rect -1049 -1588 -1015 1588
rect -791 -1588 -757 1588
rect -533 -1588 -499 1588
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
rect 499 -1588 533 1588
rect 757 -1588 791 1588
rect 1015 -1588 1049 1588
rect 1273 -1588 1307 1588
rect 1531 -1588 1565 1588
rect 1789 -1588 1823 1588
rect 2047 -1588 2081 1588
rect 2305 -1588 2339 1588
<< mvnsubdiff >>
rect -2485 1819 2485 1831
rect -2485 1785 -2377 1819
rect 2377 1785 2485 1819
rect -2485 1773 2485 1785
rect -2485 1723 -2427 1773
rect -2485 -1723 -2473 1723
rect -2439 -1723 -2427 1723
rect 2427 1723 2485 1773
rect -2485 -1773 -2427 -1723
rect 2427 -1723 2439 1723
rect 2473 -1723 2485 1723
rect 2427 -1773 2485 -1723
rect -2485 -1785 2485 -1773
rect -2485 -1819 -2377 -1785
rect 2377 -1819 2485 -1785
rect -2485 -1831 2485 -1819
<< mvnsubdiffcont >>
rect -2377 1785 2377 1819
rect -2473 -1723 -2439 1723
rect 2439 -1723 2473 1723
rect -2377 -1819 2377 -1785
<< poly >>
rect -2293 1681 -2093 1697
rect -2293 1647 -2277 1681
rect -2109 1647 -2093 1681
rect -2293 1600 -2093 1647
rect -2035 1681 -1835 1697
rect -2035 1647 -2019 1681
rect -1851 1647 -1835 1681
rect -2035 1600 -1835 1647
rect -1777 1681 -1577 1697
rect -1777 1647 -1761 1681
rect -1593 1647 -1577 1681
rect -1777 1600 -1577 1647
rect -1519 1681 -1319 1697
rect -1519 1647 -1503 1681
rect -1335 1647 -1319 1681
rect -1519 1600 -1319 1647
rect -1261 1681 -1061 1697
rect -1261 1647 -1245 1681
rect -1077 1647 -1061 1681
rect -1261 1600 -1061 1647
rect -1003 1681 -803 1697
rect -1003 1647 -987 1681
rect -819 1647 -803 1681
rect -1003 1600 -803 1647
rect -745 1681 -545 1697
rect -745 1647 -729 1681
rect -561 1647 -545 1681
rect -745 1600 -545 1647
rect -487 1681 -287 1697
rect -487 1647 -471 1681
rect -303 1647 -287 1681
rect -487 1600 -287 1647
rect -229 1681 -29 1697
rect -229 1647 -213 1681
rect -45 1647 -29 1681
rect -229 1600 -29 1647
rect 29 1681 229 1697
rect 29 1647 45 1681
rect 213 1647 229 1681
rect 29 1600 229 1647
rect 287 1681 487 1697
rect 287 1647 303 1681
rect 471 1647 487 1681
rect 287 1600 487 1647
rect 545 1681 745 1697
rect 545 1647 561 1681
rect 729 1647 745 1681
rect 545 1600 745 1647
rect 803 1681 1003 1697
rect 803 1647 819 1681
rect 987 1647 1003 1681
rect 803 1600 1003 1647
rect 1061 1681 1261 1697
rect 1061 1647 1077 1681
rect 1245 1647 1261 1681
rect 1061 1600 1261 1647
rect 1319 1681 1519 1697
rect 1319 1647 1335 1681
rect 1503 1647 1519 1681
rect 1319 1600 1519 1647
rect 1577 1681 1777 1697
rect 1577 1647 1593 1681
rect 1761 1647 1777 1681
rect 1577 1600 1777 1647
rect 1835 1681 2035 1697
rect 1835 1647 1851 1681
rect 2019 1647 2035 1681
rect 1835 1600 2035 1647
rect 2093 1681 2293 1697
rect 2093 1647 2109 1681
rect 2277 1647 2293 1681
rect 2093 1600 2293 1647
rect -2293 -1647 -2093 -1600
rect -2293 -1681 -2277 -1647
rect -2109 -1681 -2093 -1647
rect -2293 -1697 -2093 -1681
rect -2035 -1647 -1835 -1600
rect -2035 -1681 -2019 -1647
rect -1851 -1681 -1835 -1647
rect -2035 -1697 -1835 -1681
rect -1777 -1647 -1577 -1600
rect -1777 -1681 -1761 -1647
rect -1593 -1681 -1577 -1647
rect -1777 -1697 -1577 -1681
rect -1519 -1647 -1319 -1600
rect -1519 -1681 -1503 -1647
rect -1335 -1681 -1319 -1647
rect -1519 -1697 -1319 -1681
rect -1261 -1647 -1061 -1600
rect -1261 -1681 -1245 -1647
rect -1077 -1681 -1061 -1647
rect -1261 -1697 -1061 -1681
rect -1003 -1647 -803 -1600
rect -1003 -1681 -987 -1647
rect -819 -1681 -803 -1647
rect -1003 -1697 -803 -1681
rect -745 -1647 -545 -1600
rect -745 -1681 -729 -1647
rect -561 -1681 -545 -1647
rect -745 -1697 -545 -1681
rect -487 -1647 -287 -1600
rect -487 -1681 -471 -1647
rect -303 -1681 -287 -1647
rect -487 -1697 -287 -1681
rect -229 -1647 -29 -1600
rect -229 -1681 -213 -1647
rect -45 -1681 -29 -1647
rect -229 -1697 -29 -1681
rect 29 -1647 229 -1600
rect 29 -1681 45 -1647
rect 213 -1681 229 -1647
rect 29 -1697 229 -1681
rect 287 -1647 487 -1600
rect 287 -1681 303 -1647
rect 471 -1681 487 -1647
rect 287 -1697 487 -1681
rect 545 -1647 745 -1600
rect 545 -1681 561 -1647
rect 729 -1681 745 -1647
rect 545 -1697 745 -1681
rect 803 -1647 1003 -1600
rect 803 -1681 819 -1647
rect 987 -1681 1003 -1647
rect 803 -1697 1003 -1681
rect 1061 -1647 1261 -1600
rect 1061 -1681 1077 -1647
rect 1245 -1681 1261 -1647
rect 1061 -1697 1261 -1681
rect 1319 -1647 1519 -1600
rect 1319 -1681 1335 -1647
rect 1503 -1681 1519 -1647
rect 1319 -1697 1519 -1681
rect 1577 -1647 1777 -1600
rect 1577 -1681 1593 -1647
rect 1761 -1681 1777 -1647
rect 1577 -1697 1777 -1681
rect 1835 -1647 2035 -1600
rect 1835 -1681 1851 -1647
rect 2019 -1681 2035 -1647
rect 1835 -1697 2035 -1681
rect 2093 -1647 2293 -1600
rect 2093 -1681 2109 -1647
rect 2277 -1681 2293 -1647
rect 2093 -1697 2293 -1681
<< polycont >>
rect -2277 1647 -2109 1681
rect -2019 1647 -1851 1681
rect -1761 1647 -1593 1681
rect -1503 1647 -1335 1681
rect -1245 1647 -1077 1681
rect -987 1647 -819 1681
rect -729 1647 -561 1681
rect -471 1647 -303 1681
rect -213 1647 -45 1681
rect 45 1647 213 1681
rect 303 1647 471 1681
rect 561 1647 729 1681
rect 819 1647 987 1681
rect 1077 1647 1245 1681
rect 1335 1647 1503 1681
rect 1593 1647 1761 1681
rect 1851 1647 2019 1681
rect 2109 1647 2277 1681
rect -2277 -1681 -2109 -1647
rect -2019 -1681 -1851 -1647
rect -1761 -1681 -1593 -1647
rect -1503 -1681 -1335 -1647
rect -1245 -1681 -1077 -1647
rect -987 -1681 -819 -1647
rect -729 -1681 -561 -1647
rect -471 -1681 -303 -1647
rect -213 -1681 -45 -1647
rect 45 -1681 213 -1647
rect 303 -1681 471 -1647
rect 561 -1681 729 -1647
rect 819 -1681 987 -1647
rect 1077 -1681 1245 -1647
rect 1335 -1681 1503 -1647
rect 1593 -1681 1761 -1647
rect 1851 -1681 2019 -1647
rect 2109 -1681 2277 -1647
<< locali >>
rect -2473 1785 -2377 1819
rect 2377 1785 2473 1819
rect -2473 1723 -2439 1785
rect 2439 1723 2473 1785
rect -2293 1647 -2277 1681
rect -2109 1647 -2093 1681
rect -2035 1647 -2019 1681
rect -1851 1647 -1835 1681
rect -1777 1647 -1761 1681
rect -1593 1647 -1577 1681
rect -1519 1647 -1503 1681
rect -1335 1647 -1319 1681
rect -1261 1647 -1245 1681
rect -1077 1647 -1061 1681
rect -1003 1647 -987 1681
rect -819 1647 -803 1681
rect -745 1647 -729 1681
rect -561 1647 -545 1681
rect -487 1647 -471 1681
rect -303 1647 -287 1681
rect -229 1647 -213 1681
rect -45 1647 -29 1681
rect 29 1647 45 1681
rect 213 1647 229 1681
rect 287 1647 303 1681
rect 471 1647 487 1681
rect 545 1647 561 1681
rect 729 1647 745 1681
rect 803 1647 819 1681
rect 987 1647 1003 1681
rect 1061 1647 1077 1681
rect 1245 1647 1261 1681
rect 1319 1647 1335 1681
rect 1503 1647 1519 1681
rect 1577 1647 1593 1681
rect 1761 1647 1777 1681
rect 1835 1647 1851 1681
rect 2019 1647 2035 1681
rect 2093 1647 2109 1681
rect 2277 1647 2293 1681
rect -2339 1588 -2305 1604
rect -2339 -1604 -2305 -1588
rect -2081 1588 -2047 1604
rect -2081 -1604 -2047 -1588
rect -1823 1588 -1789 1604
rect -1823 -1604 -1789 -1588
rect -1565 1588 -1531 1604
rect -1565 -1604 -1531 -1588
rect -1307 1588 -1273 1604
rect -1307 -1604 -1273 -1588
rect -1049 1588 -1015 1604
rect -1049 -1604 -1015 -1588
rect -791 1588 -757 1604
rect -791 -1604 -757 -1588
rect -533 1588 -499 1604
rect -533 -1604 -499 -1588
rect -275 1588 -241 1604
rect -275 -1604 -241 -1588
rect -17 1588 17 1604
rect -17 -1604 17 -1588
rect 241 1588 275 1604
rect 241 -1604 275 -1588
rect 499 1588 533 1604
rect 499 -1604 533 -1588
rect 757 1588 791 1604
rect 757 -1604 791 -1588
rect 1015 1588 1049 1604
rect 1015 -1604 1049 -1588
rect 1273 1588 1307 1604
rect 1273 -1604 1307 -1588
rect 1531 1588 1565 1604
rect 1531 -1604 1565 -1588
rect 1789 1588 1823 1604
rect 1789 -1604 1823 -1588
rect 2047 1588 2081 1604
rect 2047 -1604 2081 -1588
rect 2305 1588 2339 1604
rect 2305 -1604 2339 -1588
rect -2293 -1681 -2277 -1647
rect -2109 -1681 -2093 -1647
rect -2035 -1681 -2019 -1647
rect -1851 -1681 -1835 -1647
rect -1777 -1681 -1761 -1647
rect -1593 -1681 -1577 -1647
rect -1519 -1681 -1503 -1647
rect -1335 -1681 -1319 -1647
rect -1261 -1681 -1245 -1647
rect -1077 -1681 -1061 -1647
rect -1003 -1681 -987 -1647
rect -819 -1681 -803 -1647
rect -745 -1681 -729 -1647
rect -561 -1681 -545 -1647
rect -487 -1681 -471 -1647
rect -303 -1681 -287 -1647
rect -229 -1681 -213 -1647
rect -45 -1681 -29 -1647
rect 29 -1681 45 -1647
rect 213 -1681 229 -1647
rect 287 -1681 303 -1647
rect 471 -1681 487 -1647
rect 545 -1681 561 -1647
rect 729 -1681 745 -1647
rect 803 -1681 819 -1647
rect 987 -1681 1003 -1647
rect 1061 -1681 1077 -1647
rect 1245 -1681 1261 -1647
rect 1319 -1681 1335 -1647
rect 1503 -1681 1519 -1647
rect 1577 -1681 1593 -1647
rect 1761 -1681 1777 -1647
rect 1835 -1681 1851 -1647
rect 2019 -1681 2035 -1647
rect 2093 -1681 2109 -1647
rect 2277 -1681 2293 -1647
rect -2473 -1785 -2439 -1723
rect 2439 -1785 2473 -1723
rect -2473 -1819 -2377 -1785
rect 2377 -1819 2473 -1785
<< viali >>
rect -2277 1647 -2109 1681
rect -2019 1647 -1851 1681
rect -1761 1647 -1593 1681
rect -1503 1647 -1335 1681
rect -1245 1647 -1077 1681
rect -987 1647 -819 1681
rect -729 1647 -561 1681
rect -471 1647 -303 1681
rect -213 1647 -45 1681
rect 45 1647 213 1681
rect 303 1647 471 1681
rect 561 1647 729 1681
rect 819 1647 987 1681
rect 1077 1647 1245 1681
rect 1335 1647 1503 1681
rect 1593 1647 1761 1681
rect 1851 1647 2019 1681
rect 2109 1647 2277 1681
rect -2339 -1588 -2305 1588
rect -2081 -1588 -2047 1588
rect -1823 -1588 -1789 1588
rect -1565 -1588 -1531 1588
rect -1307 -1588 -1273 1588
rect -1049 -1588 -1015 1588
rect -791 -1588 -757 1588
rect -533 -1588 -499 1588
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
rect 499 -1588 533 1588
rect 757 -1588 791 1588
rect 1015 -1588 1049 1588
rect 1273 -1588 1307 1588
rect 1531 -1588 1565 1588
rect 1789 -1588 1823 1588
rect 2047 -1588 2081 1588
rect 2305 -1588 2339 1588
rect -2277 -1681 -2109 -1647
rect -2019 -1681 -1851 -1647
rect -1761 -1681 -1593 -1647
rect -1503 -1681 -1335 -1647
rect -1245 -1681 -1077 -1647
rect -987 -1681 -819 -1647
rect -729 -1681 -561 -1647
rect -471 -1681 -303 -1647
rect -213 -1681 -45 -1647
rect 45 -1681 213 -1647
rect 303 -1681 471 -1647
rect 561 -1681 729 -1647
rect 819 -1681 987 -1647
rect 1077 -1681 1245 -1647
rect 1335 -1681 1503 -1647
rect 1593 -1681 1761 -1647
rect 1851 -1681 2019 -1647
rect 2109 -1681 2277 -1647
<< metal1 >>
rect -2289 1681 -2097 1687
rect -2289 1647 -2277 1681
rect -2109 1647 -2097 1681
rect -2289 1641 -2097 1647
rect -2031 1681 -1839 1687
rect -2031 1647 -2019 1681
rect -1851 1647 -1839 1681
rect -2031 1641 -1839 1647
rect -1773 1681 -1581 1687
rect -1773 1647 -1761 1681
rect -1593 1647 -1581 1681
rect -1773 1641 -1581 1647
rect -1515 1681 -1323 1687
rect -1515 1647 -1503 1681
rect -1335 1647 -1323 1681
rect -1515 1641 -1323 1647
rect -1257 1681 -1065 1687
rect -1257 1647 -1245 1681
rect -1077 1647 -1065 1681
rect -1257 1641 -1065 1647
rect -999 1681 -807 1687
rect -999 1647 -987 1681
rect -819 1647 -807 1681
rect -999 1641 -807 1647
rect -741 1681 -549 1687
rect -741 1647 -729 1681
rect -561 1647 -549 1681
rect -741 1641 -549 1647
rect -483 1681 -291 1687
rect -483 1647 -471 1681
rect -303 1647 -291 1681
rect -483 1641 -291 1647
rect -225 1681 -33 1687
rect -225 1647 -213 1681
rect -45 1647 -33 1681
rect -225 1641 -33 1647
rect 33 1681 225 1687
rect 33 1647 45 1681
rect 213 1647 225 1681
rect 33 1641 225 1647
rect 291 1681 483 1687
rect 291 1647 303 1681
rect 471 1647 483 1681
rect 291 1641 483 1647
rect 549 1681 741 1687
rect 549 1647 561 1681
rect 729 1647 741 1681
rect 549 1641 741 1647
rect 807 1681 999 1687
rect 807 1647 819 1681
rect 987 1647 999 1681
rect 807 1641 999 1647
rect 1065 1681 1257 1687
rect 1065 1647 1077 1681
rect 1245 1647 1257 1681
rect 1065 1641 1257 1647
rect 1323 1681 1515 1687
rect 1323 1647 1335 1681
rect 1503 1647 1515 1681
rect 1323 1641 1515 1647
rect 1581 1681 1773 1687
rect 1581 1647 1593 1681
rect 1761 1647 1773 1681
rect 1581 1641 1773 1647
rect 1839 1681 2031 1687
rect 1839 1647 1851 1681
rect 2019 1647 2031 1681
rect 1839 1641 2031 1647
rect 2097 1681 2289 1687
rect 2097 1647 2109 1681
rect 2277 1647 2289 1681
rect 2097 1641 2289 1647
rect -2345 1588 -2299 1600
rect -2345 -1588 -2339 1588
rect -2305 -1588 -2299 1588
rect -2345 -1600 -2299 -1588
rect -2087 1588 -2041 1600
rect -2087 -1588 -2081 1588
rect -2047 -1588 -2041 1588
rect -2087 -1600 -2041 -1588
rect -1829 1588 -1783 1600
rect -1829 -1588 -1823 1588
rect -1789 -1588 -1783 1588
rect -1829 -1600 -1783 -1588
rect -1571 1588 -1525 1600
rect -1571 -1588 -1565 1588
rect -1531 -1588 -1525 1588
rect -1571 -1600 -1525 -1588
rect -1313 1588 -1267 1600
rect -1313 -1588 -1307 1588
rect -1273 -1588 -1267 1588
rect -1313 -1600 -1267 -1588
rect -1055 1588 -1009 1600
rect -1055 -1588 -1049 1588
rect -1015 -1588 -1009 1588
rect -1055 -1600 -1009 -1588
rect -797 1588 -751 1600
rect -797 -1588 -791 1588
rect -757 -1588 -751 1588
rect -797 -1600 -751 -1588
rect -539 1588 -493 1600
rect -539 -1588 -533 1588
rect -499 -1588 -493 1588
rect -539 -1600 -493 -1588
rect -281 1588 -235 1600
rect -281 -1588 -275 1588
rect -241 -1588 -235 1588
rect -281 -1600 -235 -1588
rect -23 1588 23 1600
rect -23 -1588 -17 1588
rect 17 -1588 23 1588
rect -23 -1600 23 -1588
rect 235 1588 281 1600
rect 235 -1588 241 1588
rect 275 -1588 281 1588
rect 235 -1600 281 -1588
rect 493 1588 539 1600
rect 493 -1588 499 1588
rect 533 -1588 539 1588
rect 493 -1600 539 -1588
rect 751 1588 797 1600
rect 751 -1588 757 1588
rect 791 -1588 797 1588
rect 751 -1600 797 -1588
rect 1009 1588 1055 1600
rect 1009 -1588 1015 1588
rect 1049 -1588 1055 1588
rect 1009 -1600 1055 -1588
rect 1267 1588 1313 1600
rect 1267 -1588 1273 1588
rect 1307 -1588 1313 1588
rect 1267 -1600 1313 -1588
rect 1525 1588 1571 1600
rect 1525 -1588 1531 1588
rect 1565 -1588 1571 1588
rect 1525 -1600 1571 -1588
rect 1783 1588 1829 1600
rect 1783 -1588 1789 1588
rect 1823 -1588 1829 1588
rect 1783 -1600 1829 -1588
rect 2041 1588 2087 1600
rect 2041 -1588 2047 1588
rect 2081 -1588 2087 1588
rect 2041 -1600 2087 -1588
rect 2299 1588 2345 1600
rect 2299 -1588 2305 1588
rect 2339 -1588 2345 1588
rect 2299 -1600 2345 -1588
rect -2289 -1647 -2097 -1641
rect -2289 -1681 -2277 -1647
rect -2109 -1681 -2097 -1647
rect -2289 -1687 -2097 -1681
rect -2031 -1647 -1839 -1641
rect -2031 -1681 -2019 -1647
rect -1851 -1681 -1839 -1647
rect -2031 -1687 -1839 -1681
rect -1773 -1647 -1581 -1641
rect -1773 -1681 -1761 -1647
rect -1593 -1681 -1581 -1647
rect -1773 -1687 -1581 -1681
rect -1515 -1647 -1323 -1641
rect -1515 -1681 -1503 -1647
rect -1335 -1681 -1323 -1647
rect -1515 -1687 -1323 -1681
rect -1257 -1647 -1065 -1641
rect -1257 -1681 -1245 -1647
rect -1077 -1681 -1065 -1647
rect -1257 -1687 -1065 -1681
rect -999 -1647 -807 -1641
rect -999 -1681 -987 -1647
rect -819 -1681 -807 -1647
rect -999 -1687 -807 -1681
rect -741 -1647 -549 -1641
rect -741 -1681 -729 -1647
rect -561 -1681 -549 -1647
rect -741 -1687 -549 -1681
rect -483 -1647 -291 -1641
rect -483 -1681 -471 -1647
rect -303 -1681 -291 -1647
rect -483 -1687 -291 -1681
rect -225 -1647 -33 -1641
rect -225 -1681 -213 -1647
rect -45 -1681 -33 -1647
rect -225 -1687 -33 -1681
rect 33 -1647 225 -1641
rect 33 -1681 45 -1647
rect 213 -1681 225 -1647
rect 33 -1687 225 -1681
rect 291 -1647 483 -1641
rect 291 -1681 303 -1647
rect 471 -1681 483 -1647
rect 291 -1687 483 -1681
rect 549 -1647 741 -1641
rect 549 -1681 561 -1647
rect 729 -1681 741 -1647
rect 549 -1687 741 -1681
rect 807 -1647 999 -1641
rect 807 -1681 819 -1647
rect 987 -1681 999 -1647
rect 807 -1687 999 -1681
rect 1065 -1647 1257 -1641
rect 1065 -1681 1077 -1647
rect 1245 -1681 1257 -1647
rect 1065 -1687 1257 -1681
rect 1323 -1647 1515 -1641
rect 1323 -1681 1335 -1647
rect 1503 -1681 1515 -1647
rect 1323 -1687 1515 -1681
rect 1581 -1647 1773 -1641
rect 1581 -1681 1593 -1647
rect 1761 -1681 1773 -1647
rect 1581 -1687 1773 -1681
rect 1839 -1647 2031 -1641
rect 1839 -1681 1851 -1647
rect 2019 -1681 2031 -1647
rect 1839 -1687 2031 -1681
rect 2097 -1647 2289 -1641
rect 2097 -1681 2109 -1647
rect 2277 -1681 2289 -1647
rect 2097 -1687 2289 -1681
<< properties >>
string FIXED_BBOX -2456 -1802 2456 1802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 16 l 1 m 1 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713233716
<< nwell >>
rect -3325 -1197 3325 1197
<< mvpmos >>
rect -3067 -900 -2867 900
rect -2809 -900 -2609 900
rect -2551 -900 -2351 900
rect -2293 -900 -2093 900
rect -2035 -900 -1835 900
rect -1777 -900 -1577 900
rect -1519 -900 -1319 900
rect -1261 -900 -1061 900
rect -1003 -900 -803 900
rect -745 -900 -545 900
rect -487 -900 -287 900
rect -229 -900 -29 900
rect 29 -900 229 900
rect 287 -900 487 900
rect 545 -900 745 900
rect 803 -900 1003 900
rect 1061 -900 1261 900
rect 1319 -900 1519 900
rect 1577 -900 1777 900
rect 1835 -900 2035 900
rect 2093 -900 2293 900
rect 2351 -900 2551 900
rect 2609 -900 2809 900
rect 2867 -900 3067 900
<< mvpdiff >>
rect -3125 888 -3067 900
rect -3125 -888 -3113 888
rect -3079 -888 -3067 888
rect -3125 -900 -3067 -888
rect -2867 888 -2809 900
rect -2867 -888 -2855 888
rect -2821 -888 -2809 888
rect -2867 -900 -2809 -888
rect -2609 888 -2551 900
rect -2609 -888 -2597 888
rect -2563 -888 -2551 888
rect -2609 -900 -2551 -888
rect -2351 888 -2293 900
rect -2351 -888 -2339 888
rect -2305 -888 -2293 888
rect -2351 -900 -2293 -888
rect -2093 888 -2035 900
rect -2093 -888 -2081 888
rect -2047 -888 -2035 888
rect -2093 -900 -2035 -888
rect -1835 888 -1777 900
rect -1835 -888 -1823 888
rect -1789 -888 -1777 888
rect -1835 -900 -1777 -888
rect -1577 888 -1519 900
rect -1577 -888 -1565 888
rect -1531 -888 -1519 888
rect -1577 -900 -1519 -888
rect -1319 888 -1261 900
rect -1319 -888 -1307 888
rect -1273 -888 -1261 888
rect -1319 -900 -1261 -888
rect -1061 888 -1003 900
rect -1061 -888 -1049 888
rect -1015 -888 -1003 888
rect -1061 -900 -1003 -888
rect -803 888 -745 900
rect -803 -888 -791 888
rect -757 -888 -745 888
rect -803 -900 -745 -888
rect -545 888 -487 900
rect -545 -888 -533 888
rect -499 -888 -487 888
rect -545 -900 -487 -888
rect -287 888 -229 900
rect -287 -888 -275 888
rect -241 -888 -229 888
rect -287 -900 -229 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 229 888 287 900
rect 229 -888 241 888
rect 275 -888 287 888
rect 229 -900 287 -888
rect 487 888 545 900
rect 487 -888 499 888
rect 533 -888 545 888
rect 487 -900 545 -888
rect 745 888 803 900
rect 745 -888 757 888
rect 791 -888 803 888
rect 745 -900 803 -888
rect 1003 888 1061 900
rect 1003 -888 1015 888
rect 1049 -888 1061 888
rect 1003 -900 1061 -888
rect 1261 888 1319 900
rect 1261 -888 1273 888
rect 1307 -888 1319 888
rect 1261 -900 1319 -888
rect 1519 888 1577 900
rect 1519 -888 1531 888
rect 1565 -888 1577 888
rect 1519 -900 1577 -888
rect 1777 888 1835 900
rect 1777 -888 1789 888
rect 1823 -888 1835 888
rect 1777 -900 1835 -888
rect 2035 888 2093 900
rect 2035 -888 2047 888
rect 2081 -888 2093 888
rect 2035 -900 2093 -888
rect 2293 888 2351 900
rect 2293 -888 2305 888
rect 2339 -888 2351 888
rect 2293 -900 2351 -888
rect 2551 888 2609 900
rect 2551 -888 2563 888
rect 2597 -888 2609 888
rect 2551 -900 2609 -888
rect 2809 888 2867 900
rect 2809 -888 2821 888
rect 2855 -888 2867 888
rect 2809 -900 2867 -888
rect 3067 888 3125 900
rect 3067 -888 3079 888
rect 3113 -888 3125 888
rect 3067 -900 3125 -888
<< mvpdiffc >>
rect -3113 -888 -3079 888
rect -2855 -888 -2821 888
rect -2597 -888 -2563 888
rect -2339 -888 -2305 888
rect -2081 -888 -2047 888
rect -1823 -888 -1789 888
rect -1565 -888 -1531 888
rect -1307 -888 -1273 888
rect -1049 -888 -1015 888
rect -791 -888 -757 888
rect -533 -888 -499 888
rect -275 -888 -241 888
rect -17 -888 17 888
rect 241 -888 275 888
rect 499 -888 533 888
rect 757 -888 791 888
rect 1015 -888 1049 888
rect 1273 -888 1307 888
rect 1531 -888 1565 888
rect 1789 -888 1823 888
rect 2047 -888 2081 888
rect 2305 -888 2339 888
rect 2563 -888 2597 888
rect 2821 -888 2855 888
rect 3079 -888 3113 888
<< mvnsubdiff >>
rect -3259 1119 3259 1131
rect -3259 1085 -3151 1119
rect 3151 1085 3259 1119
rect -3259 1073 3259 1085
rect -3259 1023 -3201 1073
rect -3259 -1023 -3247 1023
rect -3213 -1023 -3201 1023
rect 3201 1023 3259 1073
rect -3259 -1073 -3201 -1023
rect 3201 -1023 3213 1023
rect 3247 -1023 3259 1023
rect 3201 -1073 3259 -1023
rect -3259 -1085 3259 -1073
rect -3259 -1119 -3151 -1085
rect 3151 -1119 3259 -1085
rect -3259 -1131 3259 -1119
<< mvnsubdiffcont >>
rect -3151 1085 3151 1119
rect -3247 -1023 -3213 1023
rect 3213 -1023 3247 1023
rect -3151 -1119 3151 -1085
<< poly >>
rect -3067 981 -2867 997
rect -3067 947 -3051 981
rect -2883 947 -2867 981
rect -3067 900 -2867 947
rect -2809 981 -2609 997
rect -2809 947 -2793 981
rect -2625 947 -2609 981
rect -2809 900 -2609 947
rect -2551 981 -2351 997
rect -2551 947 -2535 981
rect -2367 947 -2351 981
rect -2551 900 -2351 947
rect -2293 981 -2093 997
rect -2293 947 -2277 981
rect -2109 947 -2093 981
rect -2293 900 -2093 947
rect -2035 981 -1835 997
rect -2035 947 -2019 981
rect -1851 947 -1835 981
rect -2035 900 -1835 947
rect -1777 981 -1577 997
rect -1777 947 -1761 981
rect -1593 947 -1577 981
rect -1777 900 -1577 947
rect -1519 981 -1319 997
rect -1519 947 -1503 981
rect -1335 947 -1319 981
rect -1519 900 -1319 947
rect -1261 981 -1061 997
rect -1261 947 -1245 981
rect -1077 947 -1061 981
rect -1261 900 -1061 947
rect -1003 981 -803 997
rect -1003 947 -987 981
rect -819 947 -803 981
rect -1003 900 -803 947
rect -745 981 -545 997
rect -745 947 -729 981
rect -561 947 -545 981
rect -745 900 -545 947
rect -487 981 -287 997
rect -487 947 -471 981
rect -303 947 -287 981
rect -487 900 -287 947
rect -229 981 -29 997
rect -229 947 -213 981
rect -45 947 -29 981
rect -229 900 -29 947
rect 29 981 229 997
rect 29 947 45 981
rect 213 947 229 981
rect 29 900 229 947
rect 287 981 487 997
rect 287 947 303 981
rect 471 947 487 981
rect 287 900 487 947
rect 545 981 745 997
rect 545 947 561 981
rect 729 947 745 981
rect 545 900 745 947
rect 803 981 1003 997
rect 803 947 819 981
rect 987 947 1003 981
rect 803 900 1003 947
rect 1061 981 1261 997
rect 1061 947 1077 981
rect 1245 947 1261 981
rect 1061 900 1261 947
rect 1319 981 1519 997
rect 1319 947 1335 981
rect 1503 947 1519 981
rect 1319 900 1519 947
rect 1577 981 1777 997
rect 1577 947 1593 981
rect 1761 947 1777 981
rect 1577 900 1777 947
rect 1835 981 2035 997
rect 1835 947 1851 981
rect 2019 947 2035 981
rect 1835 900 2035 947
rect 2093 981 2293 997
rect 2093 947 2109 981
rect 2277 947 2293 981
rect 2093 900 2293 947
rect 2351 981 2551 997
rect 2351 947 2367 981
rect 2535 947 2551 981
rect 2351 900 2551 947
rect 2609 981 2809 997
rect 2609 947 2625 981
rect 2793 947 2809 981
rect 2609 900 2809 947
rect 2867 981 3067 997
rect 2867 947 2883 981
rect 3051 947 3067 981
rect 2867 900 3067 947
rect -3067 -947 -2867 -900
rect -3067 -981 -3051 -947
rect -2883 -981 -2867 -947
rect -3067 -997 -2867 -981
rect -2809 -947 -2609 -900
rect -2809 -981 -2793 -947
rect -2625 -981 -2609 -947
rect -2809 -997 -2609 -981
rect -2551 -947 -2351 -900
rect -2551 -981 -2535 -947
rect -2367 -981 -2351 -947
rect -2551 -997 -2351 -981
rect -2293 -947 -2093 -900
rect -2293 -981 -2277 -947
rect -2109 -981 -2093 -947
rect -2293 -997 -2093 -981
rect -2035 -947 -1835 -900
rect -2035 -981 -2019 -947
rect -1851 -981 -1835 -947
rect -2035 -997 -1835 -981
rect -1777 -947 -1577 -900
rect -1777 -981 -1761 -947
rect -1593 -981 -1577 -947
rect -1777 -997 -1577 -981
rect -1519 -947 -1319 -900
rect -1519 -981 -1503 -947
rect -1335 -981 -1319 -947
rect -1519 -997 -1319 -981
rect -1261 -947 -1061 -900
rect -1261 -981 -1245 -947
rect -1077 -981 -1061 -947
rect -1261 -997 -1061 -981
rect -1003 -947 -803 -900
rect -1003 -981 -987 -947
rect -819 -981 -803 -947
rect -1003 -997 -803 -981
rect -745 -947 -545 -900
rect -745 -981 -729 -947
rect -561 -981 -545 -947
rect -745 -997 -545 -981
rect -487 -947 -287 -900
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -487 -997 -287 -981
rect -229 -947 -29 -900
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect -229 -997 -29 -981
rect 29 -947 229 -900
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 29 -997 229 -981
rect 287 -947 487 -900
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 287 -997 487 -981
rect 545 -947 745 -900
rect 545 -981 561 -947
rect 729 -981 745 -947
rect 545 -997 745 -981
rect 803 -947 1003 -900
rect 803 -981 819 -947
rect 987 -981 1003 -947
rect 803 -997 1003 -981
rect 1061 -947 1261 -900
rect 1061 -981 1077 -947
rect 1245 -981 1261 -947
rect 1061 -997 1261 -981
rect 1319 -947 1519 -900
rect 1319 -981 1335 -947
rect 1503 -981 1519 -947
rect 1319 -997 1519 -981
rect 1577 -947 1777 -900
rect 1577 -981 1593 -947
rect 1761 -981 1777 -947
rect 1577 -997 1777 -981
rect 1835 -947 2035 -900
rect 1835 -981 1851 -947
rect 2019 -981 2035 -947
rect 1835 -997 2035 -981
rect 2093 -947 2293 -900
rect 2093 -981 2109 -947
rect 2277 -981 2293 -947
rect 2093 -997 2293 -981
rect 2351 -947 2551 -900
rect 2351 -981 2367 -947
rect 2535 -981 2551 -947
rect 2351 -997 2551 -981
rect 2609 -947 2809 -900
rect 2609 -981 2625 -947
rect 2793 -981 2809 -947
rect 2609 -997 2809 -981
rect 2867 -947 3067 -900
rect 2867 -981 2883 -947
rect 3051 -981 3067 -947
rect 2867 -997 3067 -981
<< polycont >>
rect -3051 947 -2883 981
rect -2793 947 -2625 981
rect -2535 947 -2367 981
rect -2277 947 -2109 981
rect -2019 947 -1851 981
rect -1761 947 -1593 981
rect -1503 947 -1335 981
rect -1245 947 -1077 981
rect -987 947 -819 981
rect -729 947 -561 981
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect 561 947 729 981
rect 819 947 987 981
rect 1077 947 1245 981
rect 1335 947 1503 981
rect 1593 947 1761 981
rect 1851 947 2019 981
rect 2109 947 2277 981
rect 2367 947 2535 981
rect 2625 947 2793 981
rect 2883 947 3051 981
rect -3051 -981 -2883 -947
rect -2793 -981 -2625 -947
rect -2535 -981 -2367 -947
rect -2277 -981 -2109 -947
rect -2019 -981 -1851 -947
rect -1761 -981 -1593 -947
rect -1503 -981 -1335 -947
rect -1245 -981 -1077 -947
rect -987 -981 -819 -947
rect -729 -981 -561 -947
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
rect 561 -981 729 -947
rect 819 -981 987 -947
rect 1077 -981 1245 -947
rect 1335 -981 1503 -947
rect 1593 -981 1761 -947
rect 1851 -981 2019 -947
rect 2109 -981 2277 -947
rect 2367 -981 2535 -947
rect 2625 -981 2793 -947
rect 2883 -981 3051 -947
<< locali >>
rect -3247 1085 -3151 1119
rect 3151 1085 3247 1119
rect -3247 1023 -3213 1085
rect 3213 1023 3247 1085
rect -3067 947 -3051 981
rect -2883 947 -2867 981
rect -2809 947 -2793 981
rect -2625 947 -2609 981
rect -2551 947 -2535 981
rect -2367 947 -2351 981
rect -2293 947 -2277 981
rect -2109 947 -2093 981
rect -2035 947 -2019 981
rect -1851 947 -1835 981
rect -1777 947 -1761 981
rect -1593 947 -1577 981
rect -1519 947 -1503 981
rect -1335 947 -1319 981
rect -1261 947 -1245 981
rect -1077 947 -1061 981
rect -1003 947 -987 981
rect -819 947 -803 981
rect -745 947 -729 981
rect -561 947 -545 981
rect -487 947 -471 981
rect -303 947 -287 981
rect -229 947 -213 981
rect -45 947 -29 981
rect 29 947 45 981
rect 213 947 229 981
rect 287 947 303 981
rect 471 947 487 981
rect 545 947 561 981
rect 729 947 745 981
rect 803 947 819 981
rect 987 947 1003 981
rect 1061 947 1077 981
rect 1245 947 1261 981
rect 1319 947 1335 981
rect 1503 947 1519 981
rect 1577 947 1593 981
rect 1761 947 1777 981
rect 1835 947 1851 981
rect 2019 947 2035 981
rect 2093 947 2109 981
rect 2277 947 2293 981
rect 2351 947 2367 981
rect 2535 947 2551 981
rect 2609 947 2625 981
rect 2793 947 2809 981
rect 2867 947 2883 981
rect 3051 947 3067 981
rect -3113 888 -3079 904
rect -3113 -904 -3079 -888
rect -2855 888 -2821 904
rect -2855 -904 -2821 -888
rect -2597 888 -2563 904
rect -2597 -904 -2563 -888
rect -2339 888 -2305 904
rect -2339 -904 -2305 -888
rect -2081 888 -2047 904
rect -2081 -904 -2047 -888
rect -1823 888 -1789 904
rect -1823 -904 -1789 -888
rect -1565 888 -1531 904
rect -1565 -904 -1531 -888
rect -1307 888 -1273 904
rect -1307 -904 -1273 -888
rect -1049 888 -1015 904
rect -1049 -904 -1015 -888
rect -791 888 -757 904
rect -791 -904 -757 -888
rect -533 888 -499 904
rect -533 -904 -499 -888
rect -275 888 -241 904
rect -275 -904 -241 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 241 888 275 904
rect 241 -904 275 -888
rect 499 888 533 904
rect 499 -904 533 -888
rect 757 888 791 904
rect 757 -904 791 -888
rect 1015 888 1049 904
rect 1015 -904 1049 -888
rect 1273 888 1307 904
rect 1273 -904 1307 -888
rect 1531 888 1565 904
rect 1531 -904 1565 -888
rect 1789 888 1823 904
rect 1789 -904 1823 -888
rect 2047 888 2081 904
rect 2047 -904 2081 -888
rect 2305 888 2339 904
rect 2305 -904 2339 -888
rect 2563 888 2597 904
rect 2563 -904 2597 -888
rect 2821 888 2855 904
rect 2821 -904 2855 -888
rect 3079 888 3113 904
rect 3079 -904 3113 -888
rect -3067 -981 -3051 -947
rect -2883 -981 -2867 -947
rect -2809 -981 -2793 -947
rect -2625 -981 -2609 -947
rect -2551 -981 -2535 -947
rect -2367 -981 -2351 -947
rect -2293 -981 -2277 -947
rect -2109 -981 -2093 -947
rect -2035 -981 -2019 -947
rect -1851 -981 -1835 -947
rect -1777 -981 -1761 -947
rect -1593 -981 -1577 -947
rect -1519 -981 -1503 -947
rect -1335 -981 -1319 -947
rect -1261 -981 -1245 -947
rect -1077 -981 -1061 -947
rect -1003 -981 -987 -947
rect -819 -981 -803 -947
rect -745 -981 -729 -947
rect -561 -981 -545 -947
rect -487 -981 -471 -947
rect -303 -981 -287 -947
rect -229 -981 -213 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 213 -981 229 -947
rect 287 -981 303 -947
rect 471 -981 487 -947
rect 545 -981 561 -947
rect 729 -981 745 -947
rect 803 -981 819 -947
rect 987 -981 1003 -947
rect 1061 -981 1077 -947
rect 1245 -981 1261 -947
rect 1319 -981 1335 -947
rect 1503 -981 1519 -947
rect 1577 -981 1593 -947
rect 1761 -981 1777 -947
rect 1835 -981 1851 -947
rect 2019 -981 2035 -947
rect 2093 -981 2109 -947
rect 2277 -981 2293 -947
rect 2351 -981 2367 -947
rect 2535 -981 2551 -947
rect 2609 -981 2625 -947
rect 2793 -981 2809 -947
rect 2867 -981 2883 -947
rect 3051 -981 3067 -947
rect -3247 -1085 -3213 -1023
rect 3213 -1085 3247 -1023
rect -3247 -1119 -3151 -1085
rect 3151 -1119 3247 -1085
<< viali >>
rect -3051 947 -2883 981
rect -2793 947 -2625 981
rect -2535 947 -2367 981
rect -2277 947 -2109 981
rect -2019 947 -1851 981
rect -1761 947 -1593 981
rect -1503 947 -1335 981
rect -1245 947 -1077 981
rect -987 947 -819 981
rect -729 947 -561 981
rect -471 947 -303 981
rect -213 947 -45 981
rect 45 947 213 981
rect 303 947 471 981
rect 561 947 729 981
rect 819 947 987 981
rect 1077 947 1245 981
rect 1335 947 1503 981
rect 1593 947 1761 981
rect 1851 947 2019 981
rect 2109 947 2277 981
rect 2367 947 2535 981
rect 2625 947 2793 981
rect 2883 947 3051 981
rect -3113 -888 -3079 888
rect -2855 -888 -2821 888
rect -2597 -888 -2563 888
rect -2339 -888 -2305 888
rect -2081 -888 -2047 888
rect -1823 -888 -1789 888
rect -1565 -888 -1531 888
rect -1307 -888 -1273 888
rect -1049 -888 -1015 888
rect -791 -888 -757 888
rect -533 -888 -499 888
rect -275 -888 -241 888
rect -17 -888 17 888
rect 241 -888 275 888
rect 499 -888 533 888
rect 757 -888 791 888
rect 1015 -888 1049 888
rect 1273 -888 1307 888
rect 1531 -888 1565 888
rect 1789 -888 1823 888
rect 2047 -888 2081 888
rect 2305 -888 2339 888
rect 2563 -888 2597 888
rect 2821 -888 2855 888
rect 3079 -888 3113 888
rect -3051 -981 -2883 -947
rect -2793 -981 -2625 -947
rect -2535 -981 -2367 -947
rect -2277 -981 -2109 -947
rect -2019 -981 -1851 -947
rect -1761 -981 -1593 -947
rect -1503 -981 -1335 -947
rect -1245 -981 -1077 -947
rect -987 -981 -819 -947
rect -729 -981 -561 -947
rect -471 -981 -303 -947
rect -213 -981 -45 -947
rect 45 -981 213 -947
rect 303 -981 471 -947
rect 561 -981 729 -947
rect 819 -981 987 -947
rect 1077 -981 1245 -947
rect 1335 -981 1503 -947
rect 1593 -981 1761 -947
rect 1851 -981 2019 -947
rect 2109 -981 2277 -947
rect 2367 -981 2535 -947
rect 2625 -981 2793 -947
rect 2883 -981 3051 -947
<< metal1 >>
rect -3063 981 -2871 987
rect -3063 947 -3051 981
rect -2883 947 -2871 981
rect -3063 941 -2871 947
rect -2805 981 -2613 987
rect -2805 947 -2793 981
rect -2625 947 -2613 981
rect -2805 941 -2613 947
rect -2547 981 -2355 987
rect -2547 947 -2535 981
rect -2367 947 -2355 981
rect -2547 941 -2355 947
rect -2289 981 -2097 987
rect -2289 947 -2277 981
rect -2109 947 -2097 981
rect -2289 941 -2097 947
rect -2031 981 -1839 987
rect -2031 947 -2019 981
rect -1851 947 -1839 981
rect -2031 941 -1839 947
rect -1773 981 -1581 987
rect -1773 947 -1761 981
rect -1593 947 -1581 981
rect -1773 941 -1581 947
rect -1515 981 -1323 987
rect -1515 947 -1503 981
rect -1335 947 -1323 981
rect -1515 941 -1323 947
rect -1257 981 -1065 987
rect -1257 947 -1245 981
rect -1077 947 -1065 981
rect -1257 941 -1065 947
rect -999 981 -807 987
rect -999 947 -987 981
rect -819 947 -807 981
rect -999 941 -807 947
rect -741 981 -549 987
rect -741 947 -729 981
rect -561 947 -549 981
rect -741 941 -549 947
rect -483 981 -291 987
rect -483 947 -471 981
rect -303 947 -291 981
rect -483 941 -291 947
rect -225 981 -33 987
rect -225 947 -213 981
rect -45 947 -33 981
rect -225 941 -33 947
rect 33 981 225 987
rect 33 947 45 981
rect 213 947 225 981
rect 33 941 225 947
rect 291 981 483 987
rect 291 947 303 981
rect 471 947 483 981
rect 291 941 483 947
rect 549 981 741 987
rect 549 947 561 981
rect 729 947 741 981
rect 549 941 741 947
rect 807 981 999 987
rect 807 947 819 981
rect 987 947 999 981
rect 807 941 999 947
rect 1065 981 1257 987
rect 1065 947 1077 981
rect 1245 947 1257 981
rect 1065 941 1257 947
rect 1323 981 1515 987
rect 1323 947 1335 981
rect 1503 947 1515 981
rect 1323 941 1515 947
rect 1581 981 1773 987
rect 1581 947 1593 981
rect 1761 947 1773 981
rect 1581 941 1773 947
rect 1839 981 2031 987
rect 1839 947 1851 981
rect 2019 947 2031 981
rect 1839 941 2031 947
rect 2097 981 2289 987
rect 2097 947 2109 981
rect 2277 947 2289 981
rect 2097 941 2289 947
rect 2355 981 2547 987
rect 2355 947 2367 981
rect 2535 947 2547 981
rect 2355 941 2547 947
rect 2613 981 2805 987
rect 2613 947 2625 981
rect 2793 947 2805 981
rect 2613 941 2805 947
rect 2871 981 3063 987
rect 2871 947 2883 981
rect 3051 947 3063 981
rect 2871 941 3063 947
rect -3119 888 -3073 900
rect -3119 -888 -3113 888
rect -3079 -888 -3073 888
rect -3119 -900 -3073 -888
rect -2861 888 -2815 900
rect -2861 -888 -2855 888
rect -2821 -888 -2815 888
rect -2861 -900 -2815 -888
rect -2603 888 -2557 900
rect -2603 -888 -2597 888
rect -2563 -888 -2557 888
rect -2603 -900 -2557 -888
rect -2345 888 -2299 900
rect -2345 -888 -2339 888
rect -2305 -888 -2299 888
rect -2345 -900 -2299 -888
rect -2087 888 -2041 900
rect -2087 -888 -2081 888
rect -2047 -888 -2041 888
rect -2087 -900 -2041 -888
rect -1829 888 -1783 900
rect -1829 -888 -1823 888
rect -1789 -888 -1783 888
rect -1829 -900 -1783 -888
rect -1571 888 -1525 900
rect -1571 -888 -1565 888
rect -1531 -888 -1525 888
rect -1571 -900 -1525 -888
rect -1313 888 -1267 900
rect -1313 -888 -1307 888
rect -1273 -888 -1267 888
rect -1313 -900 -1267 -888
rect -1055 888 -1009 900
rect -1055 -888 -1049 888
rect -1015 -888 -1009 888
rect -1055 -900 -1009 -888
rect -797 888 -751 900
rect -797 -888 -791 888
rect -757 -888 -751 888
rect -797 -900 -751 -888
rect -539 888 -493 900
rect -539 -888 -533 888
rect -499 -888 -493 888
rect -539 -900 -493 -888
rect -281 888 -235 900
rect -281 -888 -275 888
rect -241 -888 -235 888
rect -281 -900 -235 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 235 888 281 900
rect 235 -888 241 888
rect 275 -888 281 888
rect 235 -900 281 -888
rect 493 888 539 900
rect 493 -888 499 888
rect 533 -888 539 888
rect 493 -900 539 -888
rect 751 888 797 900
rect 751 -888 757 888
rect 791 -888 797 888
rect 751 -900 797 -888
rect 1009 888 1055 900
rect 1009 -888 1015 888
rect 1049 -888 1055 888
rect 1009 -900 1055 -888
rect 1267 888 1313 900
rect 1267 -888 1273 888
rect 1307 -888 1313 888
rect 1267 -900 1313 -888
rect 1525 888 1571 900
rect 1525 -888 1531 888
rect 1565 -888 1571 888
rect 1525 -900 1571 -888
rect 1783 888 1829 900
rect 1783 -888 1789 888
rect 1823 -888 1829 888
rect 1783 -900 1829 -888
rect 2041 888 2087 900
rect 2041 -888 2047 888
rect 2081 -888 2087 888
rect 2041 -900 2087 -888
rect 2299 888 2345 900
rect 2299 -888 2305 888
rect 2339 -888 2345 888
rect 2299 -900 2345 -888
rect 2557 888 2603 900
rect 2557 -888 2563 888
rect 2597 -888 2603 888
rect 2557 -900 2603 -888
rect 2815 888 2861 900
rect 2815 -888 2821 888
rect 2855 -888 2861 888
rect 2815 -900 2861 -888
rect 3073 888 3119 900
rect 3073 -888 3079 888
rect 3113 -888 3119 888
rect 3073 -900 3119 -888
rect -3063 -947 -2871 -941
rect -3063 -981 -3051 -947
rect -2883 -981 -2871 -947
rect -3063 -987 -2871 -981
rect -2805 -947 -2613 -941
rect -2805 -981 -2793 -947
rect -2625 -981 -2613 -947
rect -2805 -987 -2613 -981
rect -2547 -947 -2355 -941
rect -2547 -981 -2535 -947
rect -2367 -981 -2355 -947
rect -2547 -987 -2355 -981
rect -2289 -947 -2097 -941
rect -2289 -981 -2277 -947
rect -2109 -981 -2097 -947
rect -2289 -987 -2097 -981
rect -2031 -947 -1839 -941
rect -2031 -981 -2019 -947
rect -1851 -981 -1839 -947
rect -2031 -987 -1839 -981
rect -1773 -947 -1581 -941
rect -1773 -981 -1761 -947
rect -1593 -981 -1581 -947
rect -1773 -987 -1581 -981
rect -1515 -947 -1323 -941
rect -1515 -981 -1503 -947
rect -1335 -981 -1323 -947
rect -1515 -987 -1323 -981
rect -1257 -947 -1065 -941
rect -1257 -981 -1245 -947
rect -1077 -981 -1065 -947
rect -1257 -987 -1065 -981
rect -999 -947 -807 -941
rect -999 -981 -987 -947
rect -819 -981 -807 -947
rect -999 -987 -807 -981
rect -741 -947 -549 -941
rect -741 -981 -729 -947
rect -561 -981 -549 -947
rect -741 -987 -549 -981
rect -483 -947 -291 -941
rect -483 -981 -471 -947
rect -303 -981 -291 -947
rect -483 -987 -291 -981
rect -225 -947 -33 -941
rect -225 -981 -213 -947
rect -45 -981 -33 -947
rect -225 -987 -33 -981
rect 33 -947 225 -941
rect 33 -981 45 -947
rect 213 -981 225 -947
rect 33 -987 225 -981
rect 291 -947 483 -941
rect 291 -981 303 -947
rect 471 -981 483 -947
rect 291 -987 483 -981
rect 549 -947 741 -941
rect 549 -981 561 -947
rect 729 -981 741 -947
rect 549 -987 741 -981
rect 807 -947 999 -941
rect 807 -981 819 -947
rect 987 -981 999 -947
rect 807 -987 999 -981
rect 1065 -947 1257 -941
rect 1065 -981 1077 -947
rect 1245 -981 1257 -947
rect 1065 -987 1257 -981
rect 1323 -947 1515 -941
rect 1323 -981 1335 -947
rect 1503 -981 1515 -947
rect 1323 -987 1515 -981
rect 1581 -947 1773 -941
rect 1581 -981 1593 -947
rect 1761 -981 1773 -947
rect 1581 -987 1773 -981
rect 1839 -947 2031 -941
rect 1839 -981 1851 -947
rect 2019 -981 2031 -947
rect 1839 -987 2031 -981
rect 2097 -947 2289 -941
rect 2097 -981 2109 -947
rect 2277 -981 2289 -947
rect 2097 -987 2289 -981
rect 2355 -947 2547 -941
rect 2355 -981 2367 -947
rect 2535 -981 2547 -947
rect 2355 -987 2547 -981
rect 2613 -947 2805 -941
rect 2613 -981 2625 -947
rect 2793 -981 2805 -947
rect 2613 -987 2805 -981
rect 2871 -947 3063 -941
rect 2871 -981 2883 -947
rect 3051 -981 3063 -947
rect 2871 -987 3063 -981
<< properties >>
string FIXED_BBOX -3230 -1102 3230 1102
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9 l 1 m 1 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713329785
<< nwell >>
rect -3583 -897 3583 897
<< mvpmos >>
rect -3325 -600 -3125 600
rect -3067 -600 -2867 600
rect -2809 -600 -2609 600
rect -2551 -600 -2351 600
rect -2293 -600 -2093 600
rect -2035 -600 -1835 600
rect -1777 -600 -1577 600
rect -1519 -600 -1319 600
rect -1261 -600 -1061 600
rect -1003 -600 -803 600
rect -745 -600 -545 600
rect -487 -600 -287 600
rect -229 -600 -29 600
rect 29 -600 229 600
rect 287 -600 487 600
rect 545 -600 745 600
rect 803 -600 1003 600
rect 1061 -600 1261 600
rect 1319 -600 1519 600
rect 1577 -600 1777 600
rect 1835 -600 2035 600
rect 2093 -600 2293 600
rect 2351 -600 2551 600
rect 2609 -600 2809 600
rect 2867 -600 3067 600
rect 3125 -600 3325 600
<< mvpdiff >>
rect -3383 588 -3325 600
rect -3383 -588 -3371 588
rect -3337 -588 -3325 588
rect -3383 -600 -3325 -588
rect -3125 588 -3067 600
rect -3125 -588 -3113 588
rect -3079 -588 -3067 588
rect -3125 -600 -3067 -588
rect -2867 588 -2809 600
rect -2867 -588 -2855 588
rect -2821 -588 -2809 588
rect -2867 -600 -2809 -588
rect -2609 588 -2551 600
rect -2609 -588 -2597 588
rect -2563 -588 -2551 588
rect -2609 -600 -2551 -588
rect -2351 588 -2293 600
rect -2351 -588 -2339 588
rect -2305 -588 -2293 588
rect -2351 -600 -2293 -588
rect -2093 588 -2035 600
rect -2093 -588 -2081 588
rect -2047 -588 -2035 588
rect -2093 -600 -2035 -588
rect -1835 588 -1777 600
rect -1835 -588 -1823 588
rect -1789 -588 -1777 588
rect -1835 -600 -1777 -588
rect -1577 588 -1519 600
rect -1577 -588 -1565 588
rect -1531 -588 -1519 588
rect -1577 -600 -1519 -588
rect -1319 588 -1261 600
rect -1319 -588 -1307 588
rect -1273 -588 -1261 588
rect -1319 -600 -1261 -588
rect -1061 588 -1003 600
rect -1061 -588 -1049 588
rect -1015 -588 -1003 588
rect -1061 -600 -1003 -588
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -545 588 -487 600
rect -545 -588 -533 588
rect -499 -588 -487 588
rect -545 -600 -487 -588
rect -287 588 -229 600
rect -287 -588 -275 588
rect -241 -588 -229 588
rect -287 -600 -229 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 229 588 287 600
rect 229 -588 241 588
rect 275 -588 287 588
rect 229 -600 287 -588
rect 487 588 545 600
rect 487 -588 499 588
rect 533 -588 545 588
rect 487 -600 545 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
rect 1003 588 1061 600
rect 1003 -588 1015 588
rect 1049 -588 1061 588
rect 1003 -600 1061 -588
rect 1261 588 1319 600
rect 1261 -588 1273 588
rect 1307 -588 1319 588
rect 1261 -600 1319 -588
rect 1519 588 1577 600
rect 1519 -588 1531 588
rect 1565 -588 1577 588
rect 1519 -600 1577 -588
rect 1777 588 1835 600
rect 1777 -588 1789 588
rect 1823 -588 1835 588
rect 1777 -600 1835 -588
rect 2035 588 2093 600
rect 2035 -588 2047 588
rect 2081 -588 2093 588
rect 2035 -600 2093 -588
rect 2293 588 2351 600
rect 2293 -588 2305 588
rect 2339 -588 2351 588
rect 2293 -600 2351 -588
rect 2551 588 2609 600
rect 2551 -588 2563 588
rect 2597 -588 2609 588
rect 2551 -600 2609 -588
rect 2809 588 2867 600
rect 2809 -588 2821 588
rect 2855 -588 2867 588
rect 2809 -600 2867 -588
rect 3067 588 3125 600
rect 3067 -588 3079 588
rect 3113 -588 3125 588
rect 3067 -600 3125 -588
rect 3325 588 3383 600
rect 3325 -588 3337 588
rect 3371 -588 3383 588
rect 3325 -600 3383 -588
<< mvpdiffc >>
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
<< mvnsubdiff >>
rect -3517 819 3517 831
rect -3517 785 -3409 819
rect 3409 785 3517 819
rect -3517 773 3517 785
rect -3517 723 -3459 773
rect -3517 -723 -3505 723
rect -3471 -723 -3459 723
rect 3459 723 3517 773
rect -3517 -773 -3459 -723
rect 3459 -723 3471 723
rect 3505 -723 3517 723
rect 3459 -773 3517 -723
rect -3517 -785 3517 -773
rect -3517 -819 -3409 -785
rect 3409 -819 3517 -785
rect -3517 -831 3517 -819
<< mvnsubdiffcont >>
rect -3409 785 3409 819
rect -3505 -723 -3471 723
rect 3471 -723 3505 723
rect -3409 -819 3409 -785
<< poly >>
rect -3325 681 -3125 697
rect -3325 647 -3309 681
rect -3141 647 -3125 681
rect -3325 600 -3125 647
rect -3067 681 -2867 697
rect -3067 647 -3051 681
rect -2883 647 -2867 681
rect -3067 600 -2867 647
rect -2809 681 -2609 697
rect -2809 647 -2793 681
rect -2625 647 -2609 681
rect -2809 600 -2609 647
rect -2551 681 -2351 697
rect -2551 647 -2535 681
rect -2367 647 -2351 681
rect -2551 600 -2351 647
rect -2293 681 -2093 697
rect -2293 647 -2277 681
rect -2109 647 -2093 681
rect -2293 600 -2093 647
rect -2035 681 -1835 697
rect -2035 647 -2019 681
rect -1851 647 -1835 681
rect -2035 600 -1835 647
rect -1777 681 -1577 697
rect -1777 647 -1761 681
rect -1593 647 -1577 681
rect -1777 600 -1577 647
rect -1519 681 -1319 697
rect -1519 647 -1503 681
rect -1335 647 -1319 681
rect -1519 600 -1319 647
rect -1261 681 -1061 697
rect -1261 647 -1245 681
rect -1077 647 -1061 681
rect -1261 600 -1061 647
rect -1003 681 -803 697
rect -1003 647 -987 681
rect -819 647 -803 681
rect -1003 600 -803 647
rect -745 681 -545 697
rect -745 647 -729 681
rect -561 647 -545 681
rect -745 600 -545 647
rect -487 681 -287 697
rect -487 647 -471 681
rect -303 647 -287 681
rect -487 600 -287 647
rect -229 681 -29 697
rect -229 647 -213 681
rect -45 647 -29 681
rect -229 600 -29 647
rect 29 681 229 697
rect 29 647 45 681
rect 213 647 229 681
rect 29 600 229 647
rect 287 681 487 697
rect 287 647 303 681
rect 471 647 487 681
rect 287 600 487 647
rect 545 681 745 697
rect 545 647 561 681
rect 729 647 745 681
rect 545 600 745 647
rect 803 681 1003 697
rect 803 647 819 681
rect 987 647 1003 681
rect 803 600 1003 647
rect 1061 681 1261 697
rect 1061 647 1077 681
rect 1245 647 1261 681
rect 1061 600 1261 647
rect 1319 681 1519 697
rect 1319 647 1335 681
rect 1503 647 1519 681
rect 1319 600 1519 647
rect 1577 681 1777 697
rect 1577 647 1593 681
rect 1761 647 1777 681
rect 1577 600 1777 647
rect 1835 681 2035 697
rect 1835 647 1851 681
rect 2019 647 2035 681
rect 1835 600 2035 647
rect 2093 681 2293 697
rect 2093 647 2109 681
rect 2277 647 2293 681
rect 2093 600 2293 647
rect 2351 681 2551 697
rect 2351 647 2367 681
rect 2535 647 2551 681
rect 2351 600 2551 647
rect 2609 681 2809 697
rect 2609 647 2625 681
rect 2793 647 2809 681
rect 2609 600 2809 647
rect 2867 681 3067 697
rect 2867 647 2883 681
rect 3051 647 3067 681
rect 2867 600 3067 647
rect 3125 681 3325 697
rect 3125 647 3141 681
rect 3309 647 3325 681
rect 3125 600 3325 647
rect -3325 -647 -3125 -600
rect -3325 -681 -3309 -647
rect -3141 -681 -3125 -647
rect -3325 -697 -3125 -681
rect -3067 -647 -2867 -600
rect -3067 -681 -3051 -647
rect -2883 -681 -2867 -647
rect -3067 -697 -2867 -681
rect -2809 -647 -2609 -600
rect -2809 -681 -2793 -647
rect -2625 -681 -2609 -647
rect -2809 -697 -2609 -681
rect -2551 -647 -2351 -600
rect -2551 -681 -2535 -647
rect -2367 -681 -2351 -647
rect -2551 -697 -2351 -681
rect -2293 -647 -2093 -600
rect -2293 -681 -2277 -647
rect -2109 -681 -2093 -647
rect -2293 -697 -2093 -681
rect -2035 -647 -1835 -600
rect -2035 -681 -2019 -647
rect -1851 -681 -1835 -647
rect -2035 -697 -1835 -681
rect -1777 -647 -1577 -600
rect -1777 -681 -1761 -647
rect -1593 -681 -1577 -647
rect -1777 -697 -1577 -681
rect -1519 -647 -1319 -600
rect -1519 -681 -1503 -647
rect -1335 -681 -1319 -647
rect -1519 -697 -1319 -681
rect -1261 -647 -1061 -600
rect -1261 -681 -1245 -647
rect -1077 -681 -1061 -647
rect -1261 -697 -1061 -681
rect -1003 -647 -803 -600
rect -1003 -681 -987 -647
rect -819 -681 -803 -647
rect -1003 -697 -803 -681
rect -745 -647 -545 -600
rect -745 -681 -729 -647
rect -561 -681 -545 -647
rect -745 -697 -545 -681
rect -487 -647 -287 -600
rect -487 -681 -471 -647
rect -303 -681 -287 -647
rect -487 -697 -287 -681
rect -229 -647 -29 -600
rect -229 -681 -213 -647
rect -45 -681 -29 -647
rect -229 -697 -29 -681
rect 29 -647 229 -600
rect 29 -681 45 -647
rect 213 -681 229 -647
rect 29 -697 229 -681
rect 287 -647 487 -600
rect 287 -681 303 -647
rect 471 -681 487 -647
rect 287 -697 487 -681
rect 545 -647 745 -600
rect 545 -681 561 -647
rect 729 -681 745 -647
rect 545 -697 745 -681
rect 803 -647 1003 -600
rect 803 -681 819 -647
rect 987 -681 1003 -647
rect 803 -697 1003 -681
rect 1061 -647 1261 -600
rect 1061 -681 1077 -647
rect 1245 -681 1261 -647
rect 1061 -697 1261 -681
rect 1319 -647 1519 -600
rect 1319 -681 1335 -647
rect 1503 -681 1519 -647
rect 1319 -697 1519 -681
rect 1577 -647 1777 -600
rect 1577 -681 1593 -647
rect 1761 -681 1777 -647
rect 1577 -697 1777 -681
rect 1835 -647 2035 -600
rect 1835 -681 1851 -647
rect 2019 -681 2035 -647
rect 1835 -697 2035 -681
rect 2093 -647 2293 -600
rect 2093 -681 2109 -647
rect 2277 -681 2293 -647
rect 2093 -697 2293 -681
rect 2351 -647 2551 -600
rect 2351 -681 2367 -647
rect 2535 -681 2551 -647
rect 2351 -697 2551 -681
rect 2609 -647 2809 -600
rect 2609 -681 2625 -647
rect 2793 -681 2809 -647
rect 2609 -697 2809 -681
rect 2867 -647 3067 -600
rect 2867 -681 2883 -647
rect 3051 -681 3067 -647
rect 2867 -697 3067 -681
rect 3125 -647 3325 -600
rect 3125 -681 3141 -647
rect 3309 -681 3325 -647
rect 3125 -697 3325 -681
<< polycont >>
rect -3309 647 -3141 681
rect -3051 647 -2883 681
rect -2793 647 -2625 681
rect -2535 647 -2367 681
rect -2277 647 -2109 681
rect -2019 647 -1851 681
rect -1761 647 -1593 681
rect -1503 647 -1335 681
rect -1245 647 -1077 681
rect -987 647 -819 681
rect -729 647 -561 681
rect -471 647 -303 681
rect -213 647 -45 681
rect 45 647 213 681
rect 303 647 471 681
rect 561 647 729 681
rect 819 647 987 681
rect 1077 647 1245 681
rect 1335 647 1503 681
rect 1593 647 1761 681
rect 1851 647 2019 681
rect 2109 647 2277 681
rect 2367 647 2535 681
rect 2625 647 2793 681
rect 2883 647 3051 681
rect 3141 647 3309 681
rect -3309 -681 -3141 -647
rect -3051 -681 -2883 -647
rect -2793 -681 -2625 -647
rect -2535 -681 -2367 -647
rect -2277 -681 -2109 -647
rect -2019 -681 -1851 -647
rect -1761 -681 -1593 -647
rect -1503 -681 -1335 -647
rect -1245 -681 -1077 -647
rect -987 -681 -819 -647
rect -729 -681 -561 -647
rect -471 -681 -303 -647
rect -213 -681 -45 -647
rect 45 -681 213 -647
rect 303 -681 471 -647
rect 561 -681 729 -647
rect 819 -681 987 -647
rect 1077 -681 1245 -647
rect 1335 -681 1503 -647
rect 1593 -681 1761 -647
rect 1851 -681 2019 -647
rect 2109 -681 2277 -647
rect 2367 -681 2535 -647
rect 2625 -681 2793 -647
rect 2883 -681 3051 -647
rect 3141 -681 3309 -647
<< locali >>
rect -3505 785 -3409 819
rect 3409 785 3505 819
rect -3505 723 -3471 785
rect 3471 723 3505 785
rect -3325 647 -3309 681
rect -3141 647 -3125 681
rect -3067 647 -3051 681
rect -2883 647 -2867 681
rect -2809 647 -2793 681
rect -2625 647 -2609 681
rect -2551 647 -2535 681
rect -2367 647 -2351 681
rect -2293 647 -2277 681
rect -2109 647 -2093 681
rect -2035 647 -2019 681
rect -1851 647 -1835 681
rect -1777 647 -1761 681
rect -1593 647 -1577 681
rect -1519 647 -1503 681
rect -1335 647 -1319 681
rect -1261 647 -1245 681
rect -1077 647 -1061 681
rect -1003 647 -987 681
rect -819 647 -803 681
rect -745 647 -729 681
rect -561 647 -545 681
rect -487 647 -471 681
rect -303 647 -287 681
rect -229 647 -213 681
rect -45 647 -29 681
rect 29 647 45 681
rect 213 647 229 681
rect 287 647 303 681
rect 471 647 487 681
rect 545 647 561 681
rect 729 647 745 681
rect 803 647 819 681
rect 987 647 1003 681
rect 1061 647 1077 681
rect 1245 647 1261 681
rect 1319 647 1335 681
rect 1503 647 1519 681
rect 1577 647 1593 681
rect 1761 647 1777 681
rect 1835 647 1851 681
rect 2019 647 2035 681
rect 2093 647 2109 681
rect 2277 647 2293 681
rect 2351 647 2367 681
rect 2535 647 2551 681
rect 2609 647 2625 681
rect 2793 647 2809 681
rect 2867 647 2883 681
rect 3051 647 3067 681
rect 3125 647 3141 681
rect 3309 647 3325 681
rect -3371 588 -3337 604
rect -3371 -604 -3337 -588
rect -3113 588 -3079 604
rect -3113 -604 -3079 -588
rect -2855 588 -2821 604
rect -2855 -604 -2821 -588
rect -2597 588 -2563 604
rect -2597 -604 -2563 -588
rect -2339 588 -2305 604
rect -2339 -604 -2305 -588
rect -2081 588 -2047 604
rect -2081 -604 -2047 -588
rect -1823 588 -1789 604
rect -1823 -604 -1789 -588
rect -1565 588 -1531 604
rect -1565 -604 -1531 -588
rect -1307 588 -1273 604
rect -1307 -604 -1273 -588
rect -1049 588 -1015 604
rect -1049 -604 -1015 -588
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -533 588 -499 604
rect -533 -604 -499 -588
rect -275 588 -241 604
rect -275 -604 -241 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 241 588 275 604
rect 241 -604 275 -588
rect 499 588 533 604
rect 499 -604 533 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect 1015 588 1049 604
rect 1015 -604 1049 -588
rect 1273 588 1307 604
rect 1273 -604 1307 -588
rect 1531 588 1565 604
rect 1531 -604 1565 -588
rect 1789 588 1823 604
rect 1789 -604 1823 -588
rect 2047 588 2081 604
rect 2047 -604 2081 -588
rect 2305 588 2339 604
rect 2305 -604 2339 -588
rect 2563 588 2597 604
rect 2563 -604 2597 -588
rect 2821 588 2855 604
rect 2821 -604 2855 -588
rect 3079 588 3113 604
rect 3079 -604 3113 -588
rect 3337 588 3371 604
rect 3337 -604 3371 -588
rect -3325 -681 -3309 -647
rect -3141 -681 -3125 -647
rect -3067 -681 -3051 -647
rect -2883 -681 -2867 -647
rect -2809 -681 -2793 -647
rect -2625 -681 -2609 -647
rect -2551 -681 -2535 -647
rect -2367 -681 -2351 -647
rect -2293 -681 -2277 -647
rect -2109 -681 -2093 -647
rect -2035 -681 -2019 -647
rect -1851 -681 -1835 -647
rect -1777 -681 -1761 -647
rect -1593 -681 -1577 -647
rect -1519 -681 -1503 -647
rect -1335 -681 -1319 -647
rect -1261 -681 -1245 -647
rect -1077 -681 -1061 -647
rect -1003 -681 -987 -647
rect -819 -681 -803 -647
rect -745 -681 -729 -647
rect -561 -681 -545 -647
rect -487 -681 -471 -647
rect -303 -681 -287 -647
rect -229 -681 -213 -647
rect -45 -681 -29 -647
rect 29 -681 45 -647
rect 213 -681 229 -647
rect 287 -681 303 -647
rect 471 -681 487 -647
rect 545 -681 561 -647
rect 729 -681 745 -647
rect 803 -681 819 -647
rect 987 -681 1003 -647
rect 1061 -681 1077 -647
rect 1245 -681 1261 -647
rect 1319 -681 1335 -647
rect 1503 -681 1519 -647
rect 1577 -681 1593 -647
rect 1761 -681 1777 -647
rect 1835 -681 1851 -647
rect 2019 -681 2035 -647
rect 2093 -681 2109 -647
rect 2277 -681 2293 -647
rect 2351 -681 2367 -647
rect 2535 -681 2551 -647
rect 2609 -681 2625 -647
rect 2793 -681 2809 -647
rect 2867 -681 2883 -647
rect 3051 -681 3067 -647
rect 3125 -681 3141 -647
rect 3309 -681 3325 -647
rect -3505 -785 -3471 -723
rect 3471 -785 3505 -723
rect -3505 -819 -3409 -785
rect 3409 -819 3505 -785
<< viali >>
rect -3309 647 -3141 681
rect -3051 647 -2883 681
rect -2793 647 -2625 681
rect -2535 647 -2367 681
rect -2277 647 -2109 681
rect -2019 647 -1851 681
rect -1761 647 -1593 681
rect -1503 647 -1335 681
rect -1245 647 -1077 681
rect -987 647 -819 681
rect -729 647 -561 681
rect -471 647 -303 681
rect -213 647 -45 681
rect 45 647 213 681
rect 303 647 471 681
rect 561 647 729 681
rect 819 647 987 681
rect 1077 647 1245 681
rect 1335 647 1503 681
rect 1593 647 1761 681
rect 1851 647 2019 681
rect 2109 647 2277 681
rect 2367 647 2535 681
rect 2625 647 2793 681
rect 2883 647 3051 681
rect 3141 647 3309 681
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
rect -3309 -681 -3141 -647
rect -3051 -681 -2883 -647
rect -2793 -681 -2625 -647
rect -2535 -681 -2367 -647
rect -2277 -681 -2109 -647
rect -2019 -681 -1851 -647
rect -1761 -681 -1593 -647
rect -1503 -681 -1335 -647
rect -1245 -681 -1077 -647
rect -987 -681 -819 -647
rect -729 -681 -561 -647
rect -471 -681 -303 -647
rect -213 -681 -45 -647
rect 45 -681 213 -647
rect 303 -681 471 -647
rect 561 -681 729 -647
rect 819 -681 987 -647
rect 1077 -681 1245 -647
rect 1335 -681 1503 -647
rect 1593 -681 1761 -647
rect 1851 -681 2019 -647
rect 2109 -681 2277 -647
rect 2367 -681 2535 -647
rect 2625 -681 2793 -647
rect 2883 -681 3051 -647
rect 3141 -681 3309 -647
<< metal1 >>
rect -3321 681 -3129 687
rect -3321 647 -3309 681
rect -3141 647 -3129 681
rect -3321 641 -3129 647
rect -3063 681 -2871 687
rect -3063 647 -3051 681
rect -2883 647 -2871 681
rect -3063 641 -2871 647
rect -2805 681 -2613 687
rect -2805 647 -2793 681
rect -2625 647 -2613 681
rect -2805 641 -2613 647
rect -2547 681 -2355 687
rect -2547 647 -2535 681
rect -2367 647 -2355 681
rect -2547 641 -2355 647
rect -2289 681 -2097 687
rect -2289 647 -2277 681
rect -2109 647 -2097 681
rect -2289 641 -2097 647
rect -2031 681 -1839 687
rect -2031 647 -2019 681
rect -1851 647 -1839 681
rect -2031 641 -1839 647
rect -1773 681 -1581 687
rect -1773 647 -1761 681
rect -1593 647 -1581 681
rect -1773 641 -1581 647
rect -1515 681 -1323 687
rect -1515 647 -1503 681
rect -1335 647 -1323 681
rect -1515 641 -1323 647
rect -1257 681 -1065 687
rect -1257 647 -1245 681
rect -1077 647 -1065 681
rect -1257 641 -1065 647
rect -999 681 -807 687
rect -999 647 -987 681
rect -819 647 -807 681
rect -999 641 -807 647
rect -741 681 -549 687
rect -741 647 -729 681
rect -561 647 -549 681
rect -741 641 -549 647
rect -483 681 -291 687
rect -483 647 -471 681
rect -303 647 -291 681
rect -483 641 -291 647
rect -225 681 -33 687
rect -225 647 -213 681
rect -45 647 -33 681
rect -225 641 -33 647
rect 33 681 225 687
rect 33 647 45 681
rect 213 647 225 681
rect 33 641 225 647
rect 291 681 483 687
rect 291 647 303 681
rect 471 647 483 681
rect 291 641 483 647
rect 549 681 741 687
rect 549 647 561 681
rect 729 647 741 681
rect 549 641 741 647
rect 807 681 999 687
rect 807 647 819 681
rect 987 647 999 681
rect 807 641 999 647
rect 1065 681 1257 687
rect 1065 647 1077 681
rect 1245 647 1257 681
rect 1065 641 1257 647
rect 1323 681 1515 687
rect 1323 647 1335 681
rect 1503 647 1515 681
rect 1323 641 1515 647
rect 1581 681 1773 687
rect 1581 647 1593 681
rect 1761 647 1773 681
rect 1581 641 1773 647
rect 1839 681 2031 687
rect 1839 647 1851 681
rect 2019 647 2031 681
rect 1839 641 2031 647
rect 2097 681 2289 687
rect 2097 647 2109 681
rect 2277 647 2289 681
rect 2097 641 2289 647
rect 2355 681 2547 687
rect 2355 647 2367 681
rect 2535 647 2547 681
rect 2355 641 2547 647
rect 2613 681 2805 687
rect 2613 647 2625 681
rect 2793 647 2805 681
rect 2613 641 2805 647
rect 2871 681 3063 687
rect 2871 647 2883 681
rect 3051 647 3063 681
rect 2871 641 3063 647
rect 3129 681 3321 687
rect 3129 647 3141 681
rect 3309 647 3321 681
rect 3129 641 3321 647
rect -3377 588 -3331 600
rect -3377 -588 -3371 588
rect -3337 -588 -3331 588
rect -3377 -600 -3331 -588
rect -3119 588 -3073 600
rect -3119 -588 -3113 588
rect -3079 -588 -3073 588
rect -3119 -600 -3073 -588
rect -2861 588 -2815 600
rect -2861 -588 -2855 588
rect -2821 -588 -2815 588
rect -2861 -600 -2815 -588
rect -2603 588 -2557 600
rect -2603 -588 -2597 588
rect -2563 -588 -2557 588
rect -2603 -600 -2557 -588
rect -2345 588 -2299 600
rect -2345 -588 -2339 588
rect -2305 -588 -2299 588
rect -2345 -600 -2299 -588
rect -2087 588 -2041 600
rect -2087 -588 -2081 588
rect -2047 -588 -2041 588
rect -2087 -600 -2041 -588
rect -1829 588 -1783 600
rect -1829 -588 -1823 588
rect -1789 -588 -1783 588
rect -1829 -600 -1783 -588
rect -1571 588 -1525 600
rect -1571 -588 -1565 588
rect -1531 -588 -1525 588
rect -1571 -600 -1525 -588
rect -1313 588 -1267 600
rect -1313 -588 -1307 588
rect -1273 -588 -1267 588
rect -1313 -600 -1267 -588
rect -1055 588 -1009 600
rect -1055 -588 -1049 588
rect -1015 -588 -1009 588
rect -1055 -600 -1009 -588
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -539 588 -493 600
rect -539 -588 -533 588
rect -499 -588 -493 588
rect -539 -600 -493 -588
rect -281 588 -235 600
rect -281 -588 -275 588
rect -241 -588 -235 588
rect -281 -600 -235 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 235 588 281 600
rect 235 -588 241 588
rect 275 -588 281 588
rect 235 -600 281 -588
rect 493 588 539 600
rect 493 -588 499 588
rect 533 -588 539 588
rect 493 -600 539 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect 1009 588 1055 600
rect 1009 -588 1015 588
rect 1049 -588 1055 588
rect 1009 -600 1055 -588
rect 1267 588 1313 600
rect 1267 -588 1273 588
rect 1307 -588 1313 588
rect 1267 -600 1313 -588
rect 1525 588 1571 600
rect 1525 -588 1531 588
rect 1565 -588 1571 588
rect 1525 -600 1571 -588
rect 1783 588 1829 600
rect 1783 -588 1789 588
rect 1823 -588 1829 588
rect 1783 -600 1829 -588
rect 2041 588 2087 600
rect 2041 -588 2047 588
rect 2081 -588 2087 588
rect 2041 -600 2087 -588
rect 2299 588 2345 600
rect 2299 -588 2305 588
rect 2339 -588 2345 588
rect 2299 -600 2345 -588
rect 2557 588 2603 600
rect 2557 -588 2563 588
rect 2597 -588 2603 588
rect 2557 -600 2603 -588
rect 2815 588 2861 600
rect 2815 -588 2821 588
rect 2855 -588 2861 588
rect 2815 -600 2861 -588
rect 3073 588 3119 600
rect 3073 -588 3079 588
rect 3113 -588 3119 588
rect 3073 -600 3119 -588
rect 3331 588 3377 600
rect 3331 -588 3337 588
rect 3371 -588 3377 588
rect 3331 -600 3377 -588
rect -3321 -647 -3129 -641
rect -3321 -681 -3309 -647
rect -3141 -681 -3129 -647
rect -3321 -687 -3129 -681
rect -3063 -647 -2871 -641
rect -3063 -681 -3051 -647
rect -2883 -681 -2871 -647
rect -3063 -687 -2871 -681
rect -2805 -647 -2613 -641
rect -2805 -681 -2793 -647
rect -2625 -681 -2613 -647
rect -2805 -687 -2613 -681
rect -2547 -647 -2355 -641
rect -2547 -681 -2535 -647
rect -2367 -681 -2355 -647
rect -2547 -687 -2355 -681
rect -2289 -647 -2097 -641
rect -2289 -681 -2277 -647
rect -2109 -681 -2097 -647
rect -2289 -687 -2097 -681
rect -2031 -647 -1839 -641
rect -2031 -681 -2019 -647
rect -1851 -681 -1839 -647
rect -2031 -687 -1839 -681
rect -1773 -647 -1581 -641
rect -1773 -681 -1761 -647
rect -1593 -681 -1581 -647
rect -1773 -687 -1581 -681
rect -1515 -647 -1323 -641
rect -1515 -681 -1503 -647
rect -1335 -681 -1323 -647
rect -1515 -687 -1323 -681
rect -1257 -647 -1065 -641
rect -1257 -681 -1245 -647
rect -1077 -681 -1065 -647
rect -1257 -687 -1065 -681
rect -999 -647 -807 -641
rect -999 -681 -987 -647
rect -819 -681 -807 -647
rect -999 -687 -807 -681
rect -741 -647 -549 -641
rect -741 -681 -729 -647
rect -561 -681 -549 -647
rect -741 -687 -549 -681
rect -483 -647 -291 -641
rect -483 -681 -471 -647
rect -303 -681 -291 -647
rect -483 -687 -291 -681
rect -225 -647 -33 -641
rect -225 -681 -213 -647
rect -45 -681 -33 -647
rect -225 -687 -33 -681
rect 33 -647 225 -641
rect 33 -681 45 -647
rect 213 -681 225 -647
rect 33 -687 225 -681
rect 291 -647 483 -641
rect 291 -681 303 -647
rect 471 -681 483 -647
rect 291 -687 483 -681
rect 549 -647 741 -641
rect 549 -681 561 -647
rect 729 -681 741 -647
rect 549 -687 741 -681
rect 807 -647 999 -641
rect 807 -681 819 -647
rect 987 -681 999 -647
rect 807 -687 999 -681
rect 1065 -647 1257 -641
rect 1065 -681 1077 -647
rect 1245 -681 1257 -647
rect 1065 -687 1257 -681
rect 1323 -647 1515 -641
rect 1323 -681 1335 -647
rect 1503 -681 1515 -647
rect 1323 -687 1515 -681
rect 1581 -647 1773 -641
rect 1581 -681 1593 -647
rect 1761 -681 1773 -647
rect 1581 -687 1773 -681
rect 1839 -647 2031 -641
rect 1839 -681 1851 -647
rect 2019 -681 2031 -647
rect 1839 -687 2031 -681
rect 2097 -647 2289 -641
rect 2097 -681 2109 -647
rect 2277 -681 2289 -647
rect 2097 -687 2289 -681
rect 2355 -647 2547 -641
rect 2355 -681 2367 -647
rect 2535 -681 2547 -647
rect 2355 -687 2547 -681
rect 2613 -647 2805 -641
rect 2613 -681 2625 -647
rect 2793 -681 2805 -647
rect 2613 -687 2805 -681
rect 2871 -647 3063 -641
rect 2871 -681 2883 -647
rect 3051 -681 3063 -647
rect 2871 -687 3063 -681
rect 3129 -647 3321 -641
rect 3129 -681 3141 -647
rect 3309 -681 3321 -647
rect 3129 -687 3321 -681
<< properties >>
string FIXED_BBOX -3488 -802 3488 802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6 l 1 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713234246
<< nwell >>
rect -2551 -5415 2551 5415
<< mvpmos >>
rect -2293 118 -2093 5118
rect -2035 118 -1835 5118
rect -1777 118 -1577 5118
rect -1519 118 -1319 5118
rect -1261 118 -1061 5118
rect -1003 118 -803 5118
rect -745 118 -545 5118
rect -487 118 -287 5118
rect -229 118 -29 5118
rect 29 118 229 5118
rect 287 118 487 5118
rect 545 118 745 5118
rect 803 118 1003 5118
rect 1061 118 1261 5118
rect 1319 118 1519 5118
rect 1577 118 1777 5118
rect 1835 118 2035 5118
rect 2093 118 2293 5118
rect -2293 -5118 -2093 -118
rect -2035 -5118 -1835 -118
rect -1777 -5118 -1577 -118
rect -1519 -5118 -1319 -118
rect -1261 -5118 -1061 -118
rect -1003 -5118 -803 -118
rect -745 -5118 -545 -118
rect -487 -5118 -287 -118
rect -229 -5118 -29 -118
rect 29 -5118 229 -118
rect 287 -5118 487 -118
rect 545 -5118 745 -118
rect 803 -5118 1003 -118
rect 1061 -5118 1261 -118
rect 1319 -5118 1519 -118
rect 1577 -5118 1777 -118
rect 1835 -5118 2035 -118
rect 2093 -5118 2293 -118
<< mvpdiff >>
rect -2351 5106 -2293 5118
rect -2351 130 -2339 5106
rect -2305 130 -2293 5106
rect -2351 118 -2293 130
rect -2093 5106 -2035 5118
rect -2093 130 -2081 5106
rect -2047 130 -2035 5106
rect -2093 118 -2035 130
rect -1835 5106 -1777 5118
rect -1835 130 -1823 5106
rect -1789 130 -1777 5106
rect -1835 118 -1777 130
rect -1577 5106 -1519 5118
rect -1577 130 -1565 5106
rect -1531 130 -1519 5106
rect -1577 118 -1519 130
rect -1319 5106 -1261 5118
rect -1319 130 -1307 5106
rect -1273 130 -1261 5106
rect -1319 118 -1261 130
rect -1061 5106 -1003 5118
rect -1061 130 -1049 5106
rect -1015 130 -1003 5106
rect -1061 118 -1003 130
rect -803 5106 -745 5118
rect -803 130 -791 5106
rect -757 130 -745 5106
rect -803 118 -745 130
rect -545 5106 -487 5118
rect -545 130 -533 5106
rect -499 130 -487 5106
rect -545 118 -487 130
rect -287 5106 -229 5118
rect -287 130 -275 5106
rect -241 130 -229 5106
rect -287 118 -229 130
rect -29 5106 29 5118
rect -29 130 -17 5106
rect 17 130 29 5106
rect -29 118 29 130
rect 229 5106 287 5118
rect 229 130 241 5106
rect 275 130 287 5106
rect 229 118 287 130
rect 487 5106 545 5118
rect 487 130 499 5106
rect 533 130 545 5106
rect 487 118 545 130
rect 745 5106 803 5118
rect 745 130 757 5106
rect 791 130 803 5106
rect 745 118 803 130
rect 1003 5106 1061 5118
rect 1003 130 1015 5106
rect 1049 130 1061 5106
rect 1003 118 1061 130
rect 1261 5106 1319 5118
rect 1261 130 1273 5106
rect 1307 130 1319 5106
rect 1261 118 1319 130
rect 1519 5106 1577 5118
rect 1519 130 1531 5106
rect 1565 130 1577 5106
rect 1519 118 1577 130
rect 1777 5106 1835 5118
rect 1777 130 1789 5106
rect 1823 130 1835 5106
rect 1777 118 1835 130
rect 2035 5106 2093 5118
rect 2035 130 2047 5106
rect 2081 130 2093 5106
rect 2035 118 2093 130
rect 2293 5106 2351 5118
rect 2293 130 2305 5106
rect 2339 130 2351 5106
rect 2293 118 2351 130
rect -2351 -130 -2293 -118
rect -2351 -5106 -2339 -130
rect -2305 -5106 -2293 -130
rect -2351 -5118 -2293 -5106
rect -2093 -130 -2035 -118
rect -2093 -5106 -2081 -130
rect -2047 -5106 -2035 -130
rect -2093 -5118 -2035 -5106
rect -1835 -130 -1777 -118
rect -1835 -5106 -1823 -130
rect -1789 -5106 -1777 -130
rect -1835 -5118 -1777 -5106
rect -1577 -130 -1519 -118
rect -1577 -5106 -1565 -130
rect -1531 -5106 -1519 -130
rect -1577 -5118 -1519 -5106
rect -1319 -130 -1261 -118
rect -1319 -5106 -1307 -130
rect -1273 -5106 -1261 -130
rect -1319 -5118 -1261 -5106
rect -1061 -130 -1003 -118
rect -1061 -5106 -1049 -130
rect -1015 -5106 -1003 -130
rect -1061 -5118 -1003 -5106
rect -803 -130 -745 -118
rect -803 -5106 -791 -130
rect -757 -5106 -745 -130
rect -803 -5118 -745 -5106
rect -545 -130 -487 -118
rect -545 -5106 -533 -130
rect -499 -5106 -487 -130
rect -545 -5118 -487 -5106
rect -287 -130 -229 -118
rect -287 -5106 -275 -130
rect -241 -5106 -229 -130
rect -287 -5118 -229 -5106
rect -29 -130 29 -118
rect -29 -5106 -17 -130
rect 17 -5106 29 -130
rect -29 -5118 29 -5106
rect 229 -130 287 -118
rect 229 -5106 241 -130
rect 275 -5106 287 -130
rect 229 -5118 287 -5106
rect 487 -130 545 -118
rect 487 -5106 499 -130
rect 533 -5106 545 -130
rect 487 -5118 545 -5106
rect 745 -130 803 -118
rect 745 -5106 757 -130
rect 791 -5106 803 -130
rect 745 -5118 803 -5106
rect 1003 -130 1061 -118
rect 1003 -5106 1015 -130
rect 1049 -5106 1061 -130
rect 1003 -5118 1061 -5106
rect 1261 -130 1319 -118
rect 1261 -5106 1273 -130
rect 1307 -5106 1319 -130
rect 1261 -5118 1319 -5106
rect 1519 -130 1577 -118
rect 1519 -5106 1531 -130
rect 1565 -5106 1577 -130
rect 1519 -5118 1577 -5106
rect 1777 -130 1835 -118
rect 1777 -5106 1789 -130
rect 1823 -5106 1835 -130
rect 1777 -5118 1835 -5106
rect 2035 -130 2093 -118
rect 2035 -5106 2047 -130
rect 2081 -5106 2093 -130
rect 2035 -5118 2093 -5106
rect 2293 -130 2351 -118
rect 2293 -5106 2305 -130
rect 2339 -5106 2351 -130
rect 2293 -5118 2351 -5106
<< mvpdiffc >>
rect -2339 130 -2305 5106
rect -2081 130 -2047 5106
rect -1823 130 -1789 5106
rect -1565 130 -1531 5106
rect -1307 130 -1273 5106
rect -1049 130 -1015 5106
rect -791 130 -757 5106
rect -533 130 -499 5106
rect -275 130 -241 5106
rect -17 130 17 5106
rect 241 130 275 5106
rect 499 130 533 5106
rect 757 130 791 5106
rect 1015 130 1049 5106
rect 1273 130 1307 5106
rect 1531 130 1565 5106
rect 1789 130 1823 5106
rect 2047 130 2081 5106
rect 2305 130 2339 5106
rect -2339 -5106 -2305 -130
rect -2081 -5106 -2047 -130
rect -1823 -5106 -1789 -130
rect -1565 -5106 -1531 -130
rect -1307 -5106 -1273 -130
rect -1049 -5106 -1015 -130
rect -791 -5106 -757 -130
rect -533 -5106 -499 -130
rect -275 -5106 -241 -130
rect -17 -5106 17 -130
rect 241 -5106 275 -130
rect 499 -5106 533 -130
rect 757 -5106 791 -130
rect 1015 -5106 1049 -130
rect 1273 -5106 1307 -130
rect 1531 -5106 1565 -130
rect 1789 -5106 1823 -130
rect 2047 -5106 2081 -130
rect 2305 -5106 2339 -130
<< mvnsubdiff >>
rect -2485 5337 2485 5349
rect -2485 5303 -2377 5337
rect 2377 5303 2485 5337
rect -2485 5291 2485 5303
rect -2485 5241 -2427 5291
rect -2485 -5241 -2473 5241
rect -2439 -5241 -2427 5241
rect 2427 5241 2485 5291
rect -2485 -5291 -2427 -5241
rect 2427 -5241 2439 5241
rect 2473 -5241 2485 5241
rect 2427 -5291 2485 -5241
rect -2485 -5303 2485 -5291
rect -2485 -5337 -2377 -5303
rect 2377 -5337 2485 -5303
rect -2485 -5349 2485 -5337
<< mvnsubdiffcont >>
rect -2377 5303 2377 5337
rect -2473 -5241 -2439 5241
rect 2439 -5241 2473 5241
rect -2377 -5337 2377 -5303
<< poly >>
rect -2293 5199 -2093 5215
rect -2293 5165 -2277 5199
rect -2109 5165 -2093 5199
rect -2293 5118 -2093 5165
rect -2035 5199 -1835 5215
rect -2035 5165 -2019 5199
rect -1851 5165 -1835 5199
rect -2035 5118 -1835 5165
rect -1777 5199 -1577 5215
rect -1777 5165 -1761 5199
rect -1593 5165 -1577 5199
rect -1777 5118 -1577 5165
rect -1519 5199 -1319 5215
rect -1519 5165 -1503 5199
rect -1335 5165 -1319 5199
rect -1519 5118 -1319 5165
rect -1261 5199 -1061 5215
rect -1261 5165 -1245 5199
rect -1077 5165 -1061 5199
rect -1261 5118 -1061 5165
rect -1003 5199 -803 5215
rect -1003 5165 -987 5199
rect -819 5165 -803 5199
rect -1003 5118 -803 5165
rect -745 5199 -545 5215
rect -745 5165 -729 5199
rect -561 5165 -545 5199
rect -745 5118 -545 5165
rect -487 5199 -287 5215
rect -487 5165 -471 5199
rect -303 5165 -287 5199
rect -487 5118 -287 5165
rect -229 5199 -29 5215
rect -229 5165 -213 5199
rect -45 5165 -29 5199
rect -229 5118 -29 5165
rect 29 5199 229 5215
rect 29 5165 45 5199
rect 213 5165 229 5199
rect 29 5118 229 5165
rect 287 5199 487 5215
rect 287 5165 303 5199
rect 471 5165 487 5199
rect 287 5118 487 5165
rect 545 5199 745 5215
rect 545 5165 561 5199
rect 729 5165 745 5199
rect 545 5118 745 5165
rect 803 5199 1003 5215
rect 803 5165 819 5199
rect 987 5165 1003 5199
rect 803 5118 1003 5165
rect 1061 5199 1261 5215
rect 1061 5165 1077 5199
rect 1245 5165 1261 5199
rect 1061 5118 1261 5165
rect 1319 5199 1519 5215
rect 1319 5165 1335 5199
rect 1503 5165 1519 5199
rect 1319 5118 1519 5165
rect 1577 5199 1777 5215
rect 1577 5165 1593 5199
rect 1761 5165 1777 5199
rect 1577 5118 1777 5165
rect 1835 5199 2035 5215
rect 1835 5165 1851 5199
rect 2019 5165 2035 5199
rect 1835 5118 2035 5165
rect 2093 5199 2293 5215
rect 2093 5165 2109 5199
rect 2277 5165 2293 5199
rect 2093 5118 2293 5165
rect -2293 71 -2093 118
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2293 21 -2093 37
rect -2035 71 -1835 118
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 118
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 118
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 118
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 118
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 118
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 118
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 118
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 118
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 118
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 118
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 118
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect 2093 71 2293 118
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2093 21 2293 37
rect -2293 -37 -2093 -21
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2293 -118 -2093 -71
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -118 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -118 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -118 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -118 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -118 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -118 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -118 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -118 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -118 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -118 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -118 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -118 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -118 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -118 2035 -71
rect 2093 -37 2293 -21
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2093 -118 2293 -71
rect -2293 -5165 -2093 -5118
rect -2293 -5199 -2277 -5165
rect -2109 -5199 -2093 -5165
rect -2293 -5215 -2093 -5199
rect -2035 -5165 -1835 -5118
rect -2035 -5199 -2019 -5165
rect -1851 -5199 -1835 -5165
rect -2035 -5215 -1835 -5199
rect -1777 -5165 -1577 -5118
rect -1777 -5199 -1761 -5165
rect -1593 -5199 -1577 -5165
rect -1777 -5215 -1577 -5199
rect -1519 -5165 -1319 -5118
rect -1519 -5199 -1503 -5165
rect -1335 -5199 -1319 -5165
rect -1519 -5215 -1319 -5199
rect -1261 -5165 -1061 -5118
rect -1261 -5199 -1245 -5165
rect -1077 -5199 -1061 -5165
rect -1261 -5215 -1061 -5199
rect -1003 -5165 -803 -5118
rect -1003 -5199 -987 -5165
rect -819 -5199 -803 -5165
rect -1003 -5215 -803 -5199
rect -745 -5165 -545 -5118
rect -745 -5199 -729 -5165
rect -561 -5199 -545 -5165
rect -745 -5215 -545 -5199
rect -487 -5165 -287 -5118
rect -487 -5199 -471 -5165
rect -303 -5199 -287 -5165
rect -487 -5215 -287 -5199
rect -229 -5165 -29 -5118
rect -229 -5199 -213 -5165
rect -45 -5199 -29 -5165
rect -229 -5215 -29 -5199
rect 29 -5165 229 -5118
rect 29 -5199 45 -5165
rect 213 -5199 229 -5165
rect 29 -5215 229 -5199
rect 287 -5165 487 -5118
rect 287 -5199 303 -5165
rect 471 -5199 487 -5165
rect 287 -5215 487 -5199
rect 545 -5165 745 -5118
rect 545 -5199 561 -5165
rect 729 -5199 745 -5165
rect 545 -5215 745 -5199
rect 803 -5165 1003 -5118
rect 803 -5199 819 -5165
rect 987 -5199 1003 -5165
rect 803 -5215 1003 -5199
rect 1061 -5165 1261 -5118
rect 1061 -5199 1077 -5165
rect 1245 -5199 1261 -5165
rect 1061 -5215 1261 -5199
rect 1319 -5165 1519 -5118
rect 1319 -5199 1335 -5165
rect 1503 -5199 1519 -5165
rect 1319 -5215 1519 -5199
rect 1577 -5165 1777 -5118
rect 1577 -5199 1593 -5165
rect 1761 -5199 1777 -5165
rect 1577 -5215 1777 -5199
rect 1835 -5165 2035 -5118
rect 1835 -5199 1851 -5165
rect 2019 -5199 2035 -5165
rect 1835 -5215 2035 -5199
rect 2093 -5165 2293 -5118
rect 2093 -5199 2109 -5165
rect 2277 -5199 2293 -5165
rect 2093 -5215 2293 -5199
<< polycont >>
rect -2277 5165 -2109 5199
rect -2019 5165 -1851 5199
rect -1761 5165 -1593 5199
rect -1503 5165 -1335 5199
rect -1245 5165 -1077 5199
rect -987 5165 -819 5199
rect -729 5165 -561 5199
rect -471 5165 -303 5199
rect -213 5165 -45 5199
rect 45 5165 213 5199
rect 303 5165 471 5199
rect 561 5165 729 5199
rect 819 5165 987 5199
rect 1077 5165 1245 5199
rect 1335 5165 1503 5199
rect 1593 5165 1761 5199
rect 1851 5165 2019 5199
rect 2109 5165 2277 5199
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect -2277 -5199 -2109 -5165
rect -2019 -5199 -1851 -5165
rect -1761 -5199 -1593 -5165
rect -1503 -5199 -1335 -5165
rect -1245 -5199 -1077 -5165
rect -987 -5199 -819 -5165
rect -729 -5199 -561 -5165
rect -471 -5199 -303 -5165
rect -213 -5199 -45 -5165
rect 45 -5199 213 -5165
rect 303 -5199 471 -5165
rect 561 -5199 729 -5165
rect 819 -5199 987 -5165
rect 1077 -5199 1245 -5165
rect 1335 -5199 1503 -5165
rect 1593 -5199 1761 -5165
rect 1851 -5199 2019 -5165
rect 2109 -5199 2277 -5165
<< locali >>
rect -2473 5303 -2377 5337
rect 2377 5303 2473 5337
rect -2473 5241 -2439 5303
rect 2439 5241 2473 5303
rect -2293 5165 -2277 5199
rect -2109 5165 -2093 5199
rect -2035 5165 -2019 5199
rect -1851 5165 -1835 5199
rect -1777 5165 -1761 5199
rect -1593 5165 -1577 5199
rect -1519 5165 -1503 5199
rect -1335 5165 -1319 5199
rect -1261 5165 -1245 5199
rect -1077 5165 -1061 5199
rect -1003 5165 -987 5199
rect -819 5165 -803 5199
rect -745 5165 -729 5199
rect -561 5165 -545 5199
rect -487 5165 -471 5199
rect -303 5165 -287 5199
rect -229 5165 -213 5199
rect -45 5165 -29 5199
rect 29 5165 45 5199
rect 213 5165 229 5199
rect 287 5165 303 5199
rect 471 5165 487 5199
rect 545 5165 561 5199
rect 729 5165 745 5199
rect 803 5165 819 5199
rect 987 5165 1003 5199
rect 1061 5165 1077 5199
rect 1245 5165 1261 5199
rect 1319 5165 1335 5199
rect 1503 5165 1519 5199
rect 1577 5165 1593 5199
rect 1761 5165 1777 5199
rect 1835 5165 1851 5199
rect 2019 5165 2035 5199
rect 2093 5165 2109 5199
rect 2277 5165 2293 5199
rect -2339 5106 -2305 5122
rect -2339 114 -2305 130
rect -2081 5106 -2047 5122
rect -2081 114 -2047 130
rect -1823 5106 -1789 5122
rect -1823 114 -1789 130
rect -1565 5106 -1531 5122
rect -1565 114 -1531 130
rect -1307 5106 -1273 5122
rect -1307 114 -1273 130
rect -1049 5106 -1015 5122
rect -1049 114 -1015 130
rect -791 5106 -757 5122
rect -791 114 -757 130
rect -533 5106 -499 5122
rect -533 114 -499 130
rect -275 5106 -241 5122
rect -275 114 -241 130
rect -17 5106 17 5122
rect -17 114 17 130
rect 241 5106 275 5122
rect 241 114 275 130
rect 499 5106 533 5122
rect 499 114 533 130
rect 757 5106 791 5122
rect 757 114 791 130
rect 1015 5106 1049 5122
rect 1015 114 1049 130
rect 1273 5106 1307 5122
rect 1273 114 1307 130
rect 1531 5106 1565 5122
rect 1531 114 1565 130
rect 1789 5106 1823 5122
rect 1789 114 1823 130
rect 2047 5106 2081 5122
rect 2047 114 2081 130
rect 2305 5106 2339 5122
rect 2305 114 2339 130
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 2093 37 2109 71
rect 2277 37 2293 71
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect -2339 -130 -2305 -114
rect -2339 -5122 -2305 -5106
rect -2081 -130 -2047 -114
rect -2081 -5122 -2047 -5106
rect -1823 -130 -1789 -114
rect -1823 -5122 -1789 -5106
rect -1565 -130 -1531 -114
rect -1565 -5122 -1531 -5106
rect -1307 -130 -1273 -114
rect -1307 -5122 -1273 -5106
rect -1049 -130 -1015 -114
rect -1049 -5122 -1015 -5106
rect -791 -130 -757 -114
rect -791 -5122 -757 -5106
rect -533 -130 -499 -114
rect -533 -5122 -499 -5106
rect -275 -130 -241 -114
rect -275 -5122 -241 -5106
rect -17 -130 17 -114
rect -17 -5122 17 -5106
rect 241 -130 275 -114
rect 241 -5122 275 -5106
rect 499 -130 533 -114
rect 499 -5122 533 -5106
rect 757 -130 791 -114
rect 757 -5122 791 -5106
rect 1015 -130 1049 -114
rect 1015 -5122 1049 -5106
rect 1273 -130 1307 -114
rect 1273 -5122 1307 -5106
rect 1531 -130 1565 -114
rect 1531 -5122 1565 -5106
rect 1789 -130 1823 -114
rect 1789 -5122 1823 -5106
rect 2047 -130 2081 -114
rect 2047 -5122 2081 -5106
rect 2305 -130 2339 -114
rect 2305 -5122 2339 -5106
rect -2293 -5199 -2277 -5165
rect -2109 -5199 -2093 -5165
rect -2035 -5199 -2019 -5165
rect -1851 -5199 -1835 -5165
rect -1777 -5199 -1761 -5165
rect -1593 -5199 -1577 -5165
rect -1519 -5199 -1503 -5165
rect -1335 -5199 -1319 -5165
rect -1261 -5199 -1245 -5165
rect -1077 -5199 -1061 -5165
rect -1003 -5199 -987 -5165
rect -819 -5199 -803 -5165
rect -745 -5199 -729 -5165
rect -561 -5199 -545 -5165
rect -487 -5199 -471 -5165
rect -303 -5199 -287 -5165
rect -229 -5199 -213 -5165
rect -45 -5199 -29 -5165
rect 29 -5199 45 -5165
rect 213 -5199 229 -5165
rect 287 -5199 303 -5165
rect 471 -5199 487 -5165
rect 545 -5199 561 -5165
rect 729 -5199 745 -5165
rect 803 -5199 819 -5165
rect 987 -5199 1003 -5165
rect 1061 -5199 1077 -5165
rect 1245 -5199 1261 -5165
rect 1319 -5199 1335 -5165
rect 1503 -5199 1519 -5165
rect 1577 -5199 1593 -5165
rect 1761 -5199 1777 -5165
rect 1835 -5199 1851 -5165
rect 2019 -5199 2035 -5165
rect 2093 -5199 2109 -5165
rect 2277 -5199 2293 -5165
rect -2473 -5303 -2439 -5241
rect 2439 -5303 2473 -5241
rect -2473 -5337 -2377 -5303
rect 2377 -5337 2473 -5303
<< viali >>
rect -2277 5165 -2109 5199
rect -2019 5165 -1851 5199
rect -1761 5165 -1593 5199
rect -1503 5165 -1335 5199
rect -1245 5165 -1077 5199
rect -987 5165 -819 5199
rect -729 5165 -561 5199
rect -471 5165 -303 5199
rect -213 5165 -45 5199
rect 45 5165 213 5199
rect 303 5165 471 5199
rect 561 5165 729 5199
rect 819 5165 987 5199
rect 1077 5165 1245 5199
rect 1335 5165 1503 5199
rect 1593 5165 1761 5199
rect 1851 5165 2019 5199
rect 2109 5165 2277 5199
rect -2339 130 -2305 5106
rect -2081 130 -2047 5106
rect -1823 130 -1789 5106
rect -1565 130 -1531 5106
rect -1307 130 -1273 5106
rect -1049 130 -1015 5106
rect -791 130 -757 5106
rect -533 130 -499 5106
rect -275 130 -241 5106
rect -17 130 17 5106
rect 241 130 275 5106
rect 499 130 533 5106
rect 757 130 791 5106
rect 1015 130 1049 5106
rect 1273 130 1307 5106
rect 1531 130 1565 5106
rect 1789 130 1823 5106
rect 2047 130 2081 5106
rect 2305 130 2339 5106
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect -2339 -5106 -2305 -130
rect -2081 -5106 -2047 -130
rect -1823 -5106 -1789 -130
rect -1565 -5106 -1531 -130
rect -1307 -5106 -1273 -130
rect -1049 -5106 -1015 -130
rect -791 -5106 -757 -130
rect -533 -5106 -499 -130
rect -275 -5106 -241 -130
rect -17 -5106 17 -130
rect 241 -5106 275 -130
rect 499 -5106 533 -130
rect 757 -5106 791 -130
rect 1015 -5106 1049 -130
rect 1273 -5106 1307 -130
rect 1531 -5106 1565 -130
rect 1789 -5106 1823 -130
rect 2047 -5106 2081 -130
rect 2305 -5106 2339 -130
rect -2277 -5199 -2109 -5165
rect -2019 -5199 -1851 -5165
rect -1761 -5199 -1593 -5165
rect -1503 -5199 -1335 -5165
rect -1245 -5199 -1077 -5165
rect -987 -5199 -819 -5165
rect -729 -5199 -561 -5165
rect -471 -5199 -303 -5165
rect -213 -5199 -45 -5165
rect 45 -5199 213 -5165
rect 303 -5199 471 -5165
rect 561 -5199 729 -5165
rect 819 -5199 987 -5165
rect 1077 -5199 1245 -5165
rect 1335 -5199 1503 -5165
rect 1593 -5199 1761 -5165
rect 1851 -5199 2019 -5165
rect 2109 -5199 2277 -5165
<< metal1 >>
rect -2289 5199 -2097 5205
rect -2289 5165 -2277 5199
rect -2109 5165 -2097 5199
rect -2289 5159 -2097 5165
rect -2031 5199 -1839 5205
rect -2031 5165 -2019 5199
rect -1851 5165 -1839 5199
rect -2031 5159 -1839 5165
rect -1773 5199 -1581 5205
rect -1773 5165 -1761 5199
rect -1593 5165 -1581 5199
rect -1773 5159 -1581 5165
rect -1515 5199 -1323 5205
rect -1515 5165 -1503 5199
rect -1335 5165 -1323 5199
rect -1515 5159 -1323 5165
rect -1257 5199 -1065 5205
rect -1257 5165 -1245 5199
rect -1077 5165 -1065 5199
rect -1257 5159 -1065 5165
rect -999 5199 -807 5205
rect -999 5165 -987 5199
rect -819 5165 -807 5199
rect -999 5159 -807 5165
rect -741 5199 -549 5205
rect -741 5165 -729 5199
rect -561 5165 -549 5199
rect -741 5159 -549 5165
rect -483 5199 -291 5205
rect -483 5165 -471 5199
rect -303 5165 -291 5199
rect -483 5159 -291 5165
rect -225 5199 -33 5205
rect -225 5165 -213 5199
rect -45 5165 -33 5199
rect -225 5159 -33 5165
rect 33 5199 225 5205
rect 33 5165 45 5199
rect 213 5165 225 5199
rect 33 5159 225 5165
rect 291 5199 483 5205
rect 291 5165 303 5199
rect 471 5165 483 5199
rect 291 5159 483 5165
rect 549 5199 741 5205
rect 549 5165 561 5199
rect 729 5165 741 5199
rect 549 5159 741 5165
rect 807 5199 999 5205
rect 807 5165 819 5199
rect 987 5165 999 5199
rect 807 5159 999 5165
rect 1065 5199 1257 5205
rect 1065 5165 1077 5199
rect 1245 5165 1257 5199
rect 1065 5159 1257 5165
rect 1323 5199 1515 5205
rect 1323 5165 1335 5199
rect 1503 5165 1515 5199
rect 1323 5159 1515 5165
rect 1581 5199 1773 5205
rect 1581 5165 1593 5199
rect 1761 5165 1773 5199
rect 1581 5159 1773 5165
rect 1839 5199 2031 5205
rect 1839 5165 1851 5199
rect 2019 5165 2031 5199
rect 1839 5159 2031 5165
rect 2097 5199 2289 5205
rect 2097 5165 2109 5199
rect 2277 5165 2289 5199
rect 2097 5159 2289 5165
rect -2345 5106 -2299 5118
rect -2345 130 -2339 5106
rect -2305 130 -2299 5106
rect -2345 118 -2299 130
rect -2087 5106 -2041 5118
rect -2087 130 -2081 5106
rect -2047 130 -2041 5106
rect -2087 118 -2041 130
rect -1829 5106 -1783 5118
rect -1829 130 -1823 5106
rect -1789 130 -1783 5106
rect -1829 118 -1783 130
rect -1571 5106 -1525 5118
rect -1571 130 -1565 5106
rect -1531 130 -1525 5106
rect -1571 118 -1525 130
rect -1313 5106 -1267 5118
rect -1313 130 -1307 5106
rect -1273 130 -1267 5106
rect -1313 118 -1267 130
rect -1055 5106 -1009 5118
rect -1055 130 -1049 5106
rect -1015 130 -1009 5106
rect -1055 118 -1009 130
rect -797 5106 -751 5118
rect -797 130 -791 5106
rect -757 130 -751 5106
rect -797 118 -751 130
rect -539 5106 -493 5118
rect -539 130 -533 5106
rect -499 130 -493 5106
rect -539 118 -493 130
rect -281 5106 -235 5118
rect -281 130 -275 5106
rect -241 130 -235 5106
rect -281 118 -235 130
rect -23 5106 23 5118
rect -23 130 -17 5106
rect 17 130 23 5106
rect -23 118 23 130
rect 235 5106 281 5118
rect 235 130 241 5106
rect 275 130 281 5106
rect 235 118 281 130
rect 493 5106 539 5118
rect 493 130 499 5106
rect 533 130 539 5106
rect 493 118 539 130
rect 751 5106 797 5118
rect 751 130 757 5106
rect 791 130 797 5106
rect 751 118 797 130
rect 1009 5106 1055 5118
rect 1009 130 1015 5106
rect 1049 130 1055 5106
rect 1009 118 1055 130
rect 1267 5106 1313 5118
rect 1267 130 1273 5106
rect 1307 130 1313 5106
rect 1267 118 1313 130
rect 1525 5106 1571 5118
rect 1525 130 1531 5106
rect 1565 130 1571 5106
rect 1525 118 1571 130
rect 1783 5106 1829 5118
rect 1783 130 1789 5106
rect 1823 130 1829 5106
rect 1783 118 1829 130
rect 2041 5106 2087 5118
rect 2041 130 2047 5106
rect 2081 130 2087 5106
rect 2041 118 2087 130
rect 2299 5106 2345 5118
rect 2299 130 2305 5106
rect 2339 130 2345 5106
rect 2299 118 2345 130
rect -2289 71 -2097 77
rect -2289 37 -2277 71
rect -2109 37 -2097 71
rect -2289 31 -2097 37
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect 2097 71 2289 77
rect 2097 37 2109 71
rect 2277 37 2289 71
rect 2097 31 2289 37
rect -2289 -37 -2097 -31
rect -2289 -71 -2277 -37
rect -2109 -71 -2097 -37
rect -2289 -77 -2097 -71
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect 2097 -37 2289 -31
rect 2097 -71 2109 -37
rect 2277 -71 2289 -37
rect 2097 -77 2289 -71
rect -2345 -130 -2299 -118
rect -2345 -5106 -2339 -130
rect -2305 -5106 -2299 -130
rect -2345 -5118 -2299 -5106
rect -2087 -130 -2041 -118
rect -2087 -5106 -2081 -130
rect -2047 -5106 -2041 -130
rect -2087 -5118 -2041 -5106
rect -1829 -130 -1783 -118
rect -1829 -5106 -1823 -130
rect -1789 -5106 -1783 -130
rect -1829 -5118 -1783 -5106
rect -1571 -130 -1525 -118
rect -1571 -5106 -1565 -130
rect -1531 -5106 -1525 -130
rect -1571 -5118 -1525 -5106
rect -1313 -130 -1267 -118
rect -1313 -5106 -1307 -130
rect -1273 -5106 -1267 -130
rect -1313 -5118 -1267 -5106
rect -1055 -130 -1009 -118
rect -1055 -5106 -1049 -130
rect -1015 -5106 -1009 -130
rect -1055 -5118 -1009 -5106
rect -797 -130 -751 -118
rect -797 -5106 -791 -130
rect -757 -5106 -751 -130
rect -797 -5118 -751 -5106
rect -539 -130 -493 -118
rect -539 -5106 -533 -130
rect -499 -5106 -493 -130
rect -539 -5118 -493 -5106
rect -281 -130 -235 -118
rect -281 -5106 -275 -130
rect -241 -5106 -235 -130
rect -281 -5118 -235 -5106
rect -23 -130 23 -118
rect -23 -5106 -17 -130
rect 17 -5106 23 -130
rect -23 -5118 23 -5106
rect 235 -130 281 -118
rect 235 -5106 241 -130
rect 275 -5106 281 -130
rect 235 -5118 281 -5106
rect 493 -130 539 -118
rect 493 -5106 499 -130
rect 533 -5106 539 -130
rect 493 -5118 539 -5106
rect 751 -130 797 -118
rect 751 -5106 757 -130
rect 791 -5106 797 -130
rect 751 -5118 797 -5106
rect 1009 -130 1055 -118
rect 1009 -5106 1015 -130
rect 1049 -5106 1055 -130
rect 1009 -5118 1055 -5106
rect 1267 -130 1313 -118
rect 1267 -5106 1273 -130
rect 1307 -5106 1313 -130
rect 1267 -5118 1313 -5106
rect 1525 -130 1571 -118
rect 1525 -5106 1531 -130
rect 1565 -5106 1571 -130
rect 1525 -5118 1571 -5106
rect 1783 -130 1829 -118
rect 1783 -5106 1789 -130
rect 1823 -5106 1829 -130
rect 1783 -5118 1829 -5106
rect 2041 -130 2087 -118
rect 2041 -5106 2047 -130
rect 2081 -5106 2087 -130
rect 2041 -5118 2087 -5106
rect 2299 -130 2345 -118
rect 2299 -5106 2305 -130
rect 2339 -5106 2345 -130
rect 2299 -5118 2345 -5106
rect -2289 -5165 -2097 -5159
rect -2289 -5199 -2277 -5165
rect -2109 -5199 -2097 -5165
rect -2289 -5205 -2097 -5199
rect -2031 -5165 -1839 -5159
rect -2031 -5199 -2019 -5165
rect -1851 -5199 -1839 -5165
rect -2031 -5205 -1839 -5199
rect -1773 -5165 -1581 -5159
rect -1773 -5199 -1761 -5165
rect -1593 -5199 -1581 -5165
rect -1773 -5205 -1581 -5199
rect -1515 -5165 -1323 -5159
rect -1515 -5199 -1503 -5165
rect -1335 -5199 -1323 -5165
rect -1515 -5205 -1323 -5199
rect -1257 -5165 -1065 -5159
rect -1257 -5199 -1245 -5165
rect -1077 -5199 -1065 -5165
rect -1257 -5205 -1065 -5199
rect -999 -5165 -807 -5159
rect -999 -5199 -987 -5165
rect -819 -5199 -807 -5165
rect -999 -5205 -807 -5199
rect -741 -5165 -549 -5159
rect -741 -5199 -729 -5165
rect -561 -5199 -549 -5165
rect -741 -5205 -549 -5199
rect -483 -5165 -291 -5159
rect -483 -5199 -471 -5165
rect -303 -5199 -291 -5165
rect -483 -5205 -291 -5199
rect -225 -5165 -33 -5159
rect -225 -5199 -213 -5165
rect -45 -5199 -33 -5165
rect -225 -5205 -33 -5199
rect 33 -5165 225 -5159
rect 33 -5199 45 -5165
rect 213 -5199 225 -5165
rect 33 -5205 225 -5199
rect 291 -5165 483 -5159
rect 291 -5199 303 -5165
rect 471 -5199 483 -5165
rect 291 -5205 483 -5199
rect 549 -5165 741 -5159
rect 549 -5199 561 -5165
rect 729 -5199 741 -5165
rect 549 -5205 741 -5199
rect 807 -5165 999 -5159
rect 807 -5199 819 -5165
rect 987 -5199 999 -5165
rect 807 -5205 999 -5199
rect 1065 -5165 1257 -5159
rect 1065 -5199 1077 -5165
rect 1245 -5199 1257 -5165
rect 1065 -5205 1257 -5199
rect 1323 -5165 1515 -5159
rect 1323 -5199 1335 -5165
rect 1503 -5199 1515 -5165
rect 1323 -5205 1515 -5199
rect 1581 -5165 1773 -5159
rect 1581 -5199 1593 -5165
rect 1761 -5199 1773 -5165
rect 1581 -5205 1773 -5199
rect 1839 -5165 2031 -5159
rect 1839 -5199 1851 -5165
rect 2019 -5199 2031 -5165
rect 1839 -5205 2031 -5199
rect 2097 -5165 2289 -5159
rect 2097 -5199 2109 -5165
rect 2277 -5199 2289 -5165
rect 2097 -5205 2289 -5199
<< properties >>
string FIXED_BBOX -2456 -5320 2456 5320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 25 l 1 m 2 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

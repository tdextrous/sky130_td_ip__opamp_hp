magic
tech sky130A
magscale 1 2
timestamp 1713394428
<< nwell >>
rect -3583 -897 3583 897
<< mvpmos >>
rect -3325 -600 -3125 600
rect -3067 -600 -2867 600
rect -2809 -600 -2609 600
rect -2551 -600 -2351 600
rect -2293 -600 -2093 600
rect -2035 -600 -1835 600
rect -1777 -600 -1577 600
rect -1519 -600 -1319 600
rect -1261 -600 -1061 600
rect -1003 -600 -803 600
rect -745 -600 -545 600
rect -487 -600 -287 600
rect -229 -600 -29 600
rect 29 -600 229 600
rect 287 -600 487 600
rect 545 -600 745 600
rect 803 -600 1003 600
rect 1061 -600 1261 600
rect 1319 -600 1519 600
rect 1577 -600 1777 600
rect 1835 -600 2035 600
rect 2093 -600 2293 600
rect 2351 -600 2551 600
rect 2609 -600 2809 600
rect 2867 -600 3067 600
rect 3125 -600 3325 600
<< mvpdiff >>
rect -3383 588 -3325 600
rect -3383 -588 -3371 588
rect -3337 -588 -3325 588
rect -3383 -600 -3325 -588
rect -3125 588 -3067 600
rect -3125 -588 -3113 588
rect -3079 -588 -3067 588
rect -3125 -600 -3067 -588
rect -2867 588 -2809 600
rect -2867 -588 -2855 588
rect -2821 -588 -2809 588
rect -2867 -600 -2809 -588
rect -2609 588 -2551 600
rect -2609 -588 -2597 588
rect -2563 -588 -2551 588
rect -2609 -600 -2551 -588
rect -2351 588 -2293 600
rect -2351 -588 -2339 588
rect -2305 -588 -2293 588
rect -2351 -600 -2293 -588
rect -2093 588 -2035 600
rect -2093 -588 -2081 588
rect -2047 -588 -2035 588
rect -2093 -600 -2035 -588
rect -1835 588 -1777 600
rect -1835 -588 -1823 588
rect -1789 -588 -1777 588
rect -1835 -600 -1777 -588
rect -1577 588 -1519 600
rect -1577 -588 -1565 588
rect -1531 -588 -1519 588
rect -1577 -600 -1519 -588
rect -1319 588 -1261 600
rect -1319 -588 -1307 588
rect -1273 -588 -1261 588
rect -1319 -600 -1261 -588
rect -1061 588 -1003 600
rect -1061 -588 -1049 588
rect -1015 -588 -1003 588
rect -1061 -600 -1003 -588
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -545 588 -487 600
rect -545 -588 -533 588
rect -499 -588 -487 588
rect -545 -600 -487 -588
rect -287 588 -229 600
rect -287 -588 -275 588
rect -241 -588 -229 588
rect -287 -600 -229 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 229 588 287 600
rect 229 -588 241 588
rect 275 -588 287 588
rect 229 -600 287 -588
rect 487 588 545 600
rect 487 -588 499 588
rect 533 -588 545 588
rect 487 -600 545 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
rect 1003 588 1061 600
rect 1003 -588 1015 588
rect 1049 -588 1061 588
rect 1003 -600 1061 -588
rect 1261 588 1319 600
rect 1261 -588 1273 588
rect 1307 -588 1319 588
rect 1261 -600 1319 -588
rect 1519 588 1577 600
rect 1519 -588 1531 588
rect 1565 -588 1577 588
rect 1519 -600 1577 -588
rect 1777 588 1835 600
rect 1777 -588 1789 588
rect 1823 -588 1835 588
rect 1777 -600 1835 -588
rect 2035 588 2093 600
rect 2035 -588 2047 588
rect 2081 -588 2093 588
rect 2035 -600 2093 -588
rect 2293 588 2351 600
rect 2293 -588 2305 588
rect 2339 -588 2351 588
rect 2293 -600 2351 -588
rect 2551 588 2609 600
rect 2551 -588 2563 588
rect 2597 -588 2609 588
rect 2551 -600 2609 -588
rect 2809 588 2867 600
rect 2809 -588 2821 588
rect 2855 -588 2867 588
rect 2809 -600 2867 -588
rect 3067 588 3125 600
rect 3067 -588 3079 588
rect 3113 -588 3125 588
rect 3067 -600 3125 -588
rect 3325 588 3383 600
rect 3325 -588 3337 588
rect 3371 -588 3383 588
rect 3325 -600 3383 -588
<< mvpdiffc >>
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
<< mvnsubdiff >>
rect -3517 819 3517 831
rect -3517 785 -3409 819
rect 3409 785 3517 819
rect -3517 773 3517 785
rect -3517 723 -3459 773
rect -3517 -723 -3505 723
rect -3471 -723 -3459 723
rect 3459 723 3517 773
rect -3517 -773 -3459 -723
rect 3459 -723 3471 723
rect 3505 -723 3517 723
rect 3459 -773 3517 -723
rect -3517 -785 3517 -773
rect -3517 -819 -3409 -785
rect 3409 -819 3517 -785
rect -3517 -831 3517 -819
<< mvnsubdiffcont >>
rect -3409 785 3409 819
rect -3505 -723 -3471 723
rect 3471 -723 3505 723
rect -3409 -819 3409 -785
<< poly >>
rect -3291 681 -3159 697
rect -3291 664 -3275 681
rect -3325 647 -3275 664
rect -3175 664 -3159 681
rect -3033 681 -2901 697
rect -3033 664 -3017 681
rect -3175 647 -3125 664
rect -3325 600 -3125 647
rect -3067 647 -3017 664
rect -2917 664 -2901 681
rect -2775 681 -2643 697
rect -2775 664 -2759 681
rect -2917 647 -2867 664
rect -3067 600 -2867 647
rect -2809 647 -2759 664
rect -2659 664 -2643 681
rect -2517 681 -2385 697
rect -2517 664 -2501 681
rect -2659 647 -2609 664
rect -2809 600 -2609 647
rect -2551 647 -2501 664
rect -2401 664 -2385 681
rect -2259 681 -2127 697
rect -2259 664 -2243 681
rect -2401 647 -2351 664
rect -2551 600 -2351 647
rect -2293 647 -2243 664
rect -2143 664 -2127 681
rect -2001 681 -1869 697
rect -2001 664 -1985 681
rect -2143 647 -2093 664
rect -2293 600 -2093 647
rect -2035 647 -1985 664
rect -1885 664 -1869 681
rect -1743 681 -1611 697
rect -1743 664 -1727 681
rect -1885 647 -1835 664
rect -2035 600 -1835 647
rect -1777 647 -1727 664
rect -1627 664 -1611 681
rect -1485 681 -1353 697
rect -1485 664 -1469 681
rect -1627 647 -1577 664
rect -1777 600 -1577 647
rect -1519 647 -1469 664
rect -1369 664 -1353 681
rect -1227 681 -1095 697
rect -1227 664 -1211 681
rect -1369 647 -1319 664
rect -1519 600 -1319 647
rect -1261 647 -1211 664
rect -1111 664 -1095 681
rect -969 681 -837 697
rect -969 664 -953 681
rect -1111 647 -1061 664
rect -1261 600 -1061 647
rect -1003 647 -953 664
rect -853 664 -837 681
rect -711 681 -579 697
rect -711 664 -695 681
rect -853 647 -803 664
rect -1003 600 -803 647
rect -745 647 -695 664
rect -595 664 -579 681
rect -453 681 -321 697
rect -453 664 -437 681
rect -595 647 -545 664
rect -745 600 -545 647
rect -487 647 -437 664
rect -337 664 -321 681
rect -195 681 -63 697
rect -195 664 -179 681
rect -337 647 -287 664
rect -487 600 -287 647
rect -229 647 -179 664
rect -79 664 -63 681
rect 63 681 195 697
rect 63 664 79 681
rect -79 647 -29 664
rect -229 600 -29 647
rect 29 647 79 664
rect 179 664 195 681
rect 321 681 453 697
rect 321 664 337 681
rect 179 647 229 664
rect 29 600 229 647
rect 287 647 337 664
rect 437 664 453 681
rect 579 681 711 697
rect 579 664 595 681
rect 437 647 487 664
rect 287 600 487 647
rect 545 647 595 664
rect 695 664 711 681
rect 837 681 969 697
rect 837 664 853 681
rect 695 647 745 664
rect 545 600 745 647
rect 803 647 853 664
rect 953 664 969 681
rect 1095 681 1227 697
rect 1095 664 1111 681
rect 953 647 1003 664
rect 803 600 1003 647
rect 1061 647 1111 664
rect 1211 664 1227 681
rect 1353 681 1485 697
rect 1353 664 1369 681
rect 1211 647 1261 664
rect 1061 600 1261 647
rect 1319 647 1369 664
rect 1469 664 1485 681
rect 1611 681 1743 697
rect 1611 664 1627 681
rect 1469 647 1519 664
rect 1319 600 1519 647
rect 1577 647 1627 664
rect 1727 664 1743 681
rect 1869 681 2001 697
rect 1869 664 1885 681
rect 1727 647 1777 664
rect 1577 600 1777 647
rect 1835 647 1885 664
rect 1985 664 2001 681
rect 2127 681 2259 697
rect 2127 664 2143 681
rect 1985 647 2035 664
rect 1835 600 2035 647
rect 2093 647 2143 664
rect 2243 664 2259 681
rect 2385 681 2517 697
rect 2385 664 2401 681
rect 2243 647 2293 664
rect 2093 600 2293 647
rect 2351 647 2401 664
rect 2501 664 2517 681
rect 2643 681 2775 697
rect 2643 664 2659 681
rect 2501 647 2551 664
rect 2351 600 2551 647
rect 2609 647 2659 664
rect 2759 664 2775 681
rect 2901 681 3033 697
rect 2901 664 2917 681
rect 2759 647 2809 664
rect 2609 600 2809 647
rect 2867 647 2917 664
rect 3017 664 3033 681
rect 3159 681 3291 697
rect 3159 664 3175 681
rect 3017 647 3067 664
rect 2867 600 3067 647
rect 3125 647 3175 664
rect 3275 664 3291 681
rect 3275 647 3325 664
rect 3125 600 3325 647
rect -3325 -647 -3125 -600
rect -3325 -664 -3275 -647
rect -3291 -681 -3275 -664
rect -3175 -664 -3125 -647
rect -3067 -647 -2867 -600
rect -3067 -664 -3017 -647
rect -3175 -681 -3159 -664
rect -3291 -697 -3159 -681
rect -3033 -681 -3017 -664
rect -2917 -664 -2867 -647
rect -2809 -647 -2609 -600
rect -2809 -664 -2759 -647
rect -2917 -681 -2901 -664
rect -3033 -697 -2901 -681
rect -2775 -681 -2759 -664
rect -2659 -664 -2609 -647
rect -2551 -647 -2351 -600
rect -2551 -664 -2501 -647
rect -2659 -681 -2643 -664
rect -2775 -697 -2643 -681
rect -2517 -681 -2501 -664
rect -2401 -664 -2351 -647
rect -2293 -647 -2093 -600
rect -2293 -664 -2243 -647
rect -2401 -681 -2385 -664
rect -2517 -697 -2385 -681
rect -2259 -681 -2243 -664
rect -2143 -664 -2093 -647
rect -2035 -647 -1835 -600
rect -2035 -664 -1985 -647
rect -2143 -681 -2127 -664
rect -2259 -697 -2127 -681
rect -2001 -681 -1985 -664
rect -1885 -664 -1835 -647
rect -1777 -647 -1577 -600
rect -1777 -664 -1727 -647
rect -1885 -681 -1869 -664
rect -2001 -697 -1869 -681
rect -1743 -681 -1727 -664
rect -1627 -664 -1577 -647
rect -1519 -647 -1319 -600
rect -1519 -664 -1469 -647
rect -1627 -681 -1611 -664
rect -1743 -697 -1611 -681
rect -1485 -681 -1469 -664
rect -1369 -664 -1319 -647
rect -1261 -647 -1061 -600
rect -1261 -664 -1211 -647
rect -1369 -681 -1353 -664
rect -1485 -697 -1353 -681
rect -1227 -681 -1211 -664
rect -1111 -664 -1061 -647
rect -1003 -647 -803 -600
rect -1003 -664 -953 -647
rect -1111 -681 -1095 -664
rect -1227 -697 -1095 -681
rect -969 -681 -953 -664
rect -853 -664 -803 -647
rect -745 -647 -545 -600
rect -745 -664 -695 -647
rect -853 -681 -837 -664
rect -969 -697 -837 -681
rect -711 -681 -695 -664
rect -595 -664 -545 -647
rect -487 -647 -287 -600
rect -487 -664 -437 -647
rect -595 -681 -579 -664
rect -711 -697 -579 -681
rect -453 -681 -437 -664
rect -337 -664 -287 -647
rect -229 -647 -29 -600
rect -229 -664 -179 -647
rect -337 -681 -321 -664
rect -453 -697 -321 -681
rect -195 -681 -179 -664
rect -79 -664 -29 -647
rect 29 -647 229 -600
rect 29 -664 79 -647
rect -79 -681 -63 -664
rect -195 -697 -63 -681
rect 63 -681 79 -664
rect 179 -664 229 -647
rect 287 -647 487 -600
rect 287 -664 337 -647
rect 179 -681 195 -664
rect 63 -697 195 -681
rect 321 -681 337 -664
rect 437 -664 487 -647
rect 545 -647 745 -600
rect 545 -664 595 -647
rect 437 -681 453 -664
rect 321 -697 453 -681
rect 579 -681 595 -664
rect 695 -664 745 -647
rect 803 -647 1003 -600
rect 803 -664 853 -647
rect 695 -681 711 -664
rect 579 -697 711 -681
rect 837 -681 853 -664
rect 953 -664 1003 -647
rect 1061 -647 1261 -600
rect 1061 -664 1111 -647
rect 953 -681 969 -664
rect 837 -697 969 -681
rect 1095 -681 1111 -664
rect 1211 -664 1261 -647
rect 1319 -647 1519 -600
rect 1319 -664 1369 -647
rect 1211 -681 1227 -664
rect 1095 -697 1227 -681
rect 1353 -681 1369 -664
rect 1469 -664 1519 -647
rect 1577 -647 1777 -600
rect 1577 -664 1627 -647
rect 1469 -681 1485 -664
rect 1353 -697 1485 -681
rect 1611 -681 1627 -664
rect 1727 -664 1777 -647
rect 1835 -647 2035 -600
rect 1835 -664 1885 -647
rect 1727 -681 1743 -664
rect 1611 -697 1743 -681
rect 1869 -681 1885 -664
rect 1985 -664 2035 -647
rect 2093 -647 2293 -600
rect 2093 -664 2143 -647
rect 1985 -681 2001 -664
rect 1869 -697 2001 -681
rect 2127 -681 2143 -664
rect 2243 -664 2293 -647
rect 2351 -647 2551 -600
rect 2351 -664 2401 -647
rect 2243 -681 2259 -664
rect 2127 -697 2259 -681
rect 2385 -681 2401 -664
rect 2501 -664 2551 -647
rect 2609 -647 2809 -600
rect 2609 -664 2659 -647
rect 2501 -681 2517 -664
rect 2385 -697 2517 -681
rect 2643 -681 2659 -664
rect 2759 -664 2809 -647
rect 2867 -647 3067 -600
rect 2867 -664 2917 -647
rect 2759 -681 2775 -664
rect 2643 -697 2775 -681
rect 2901 -681 2917 -664
rect 3017 -664 3067 -647
rect 3125 -647 3325 -600
rect 3125 -664 3175 -647
rect 3017 -681 3033 -664
rect 2901 -697 3033 -681
rect 3159 -681 3175 -664
rect 3275 -664 3325 -647
rect 3275 -681 3291 -664
rect 3159 -697 3291 -681
<< polycont >>
rect -3275 647 -3175 681
rect -3017 647 -2917 681
rect -2759 647 -2659 681
rect -2501 647 -2401 681
rect -2243 647 -2143 681
rect -1985 647 -1885 681
rect -1727 647 -1627 681
rect -1469 647 -1369 681
rect -1211 647 -1111 681
rect -953 647 -853 681
rect -695 647 -595 681
rect -437 647 -337 681
rect -179 647 -79 681
rect 79 647 179 681
rect 337 647 437 681
rect 595 647 695 681
rect 853 647 953 681
rect 1111 647 1211 681
rect 1369 647 1469 681
rect 1627 647 1727 681
rect 1885 647 1985 681
rect 2143 647 2243 681
rect 2401 647 2501 681
rect 2659 647 2759 681
rect 2917 647 3017 681
rect 3175 647 3275 681
rect -3275 -681 -3175 -647
rect -3017 -681 -2917 -647
rect -2759 -681 -2659 -647
rect -2501 -681 -2401 -647
rect -2243 -681 -2143 -647
rect -1985 -681 -1885 -647
rect -1727 -681 -1627 -647
rect -1469 -681 -1369 -647
rect -1211 -681 -1111 -647
rect -953 -681 -853 -647
rect -695 -681 -595 -647
rect -437 -681 -337 -647
rect -179 -681 -79 -647
rect 79 -681 179 -647
rect 337 -681 437 -647
rect 595 -681 695 -647
rect 853 -681 953 -647
rect 1111 -681 1211 -647
rect 1369 -681 1469 -647
rect 1627 -681 1727 -647
rect 1885 -681 1985 -647
rect 2143 -681 2243 -647
rect 2401 -681 2501 -647
rect 2659 -681 2759 -647
rect 2917 -681 3017 -647
rect 3175 -681 3275 -647
<< locali >>
rect -3505 785 -3409 819
rect 3409 785 3505 819
rect -3505 723 -3471 785
rect 3471 723 3505 785
rect -3291 647 -3275 681
rect -3175 647 -3159 681
rect -3033 647 -3017 681
rect -2917 647 -2901 681
rect -2775 647 -2759 681
rect -2659 647 -2643 681
rect -2517 647 -2501 681
rect -2401 647 -2385 681
rect -2259 647 -2243 681
rect -2143 647 -2127 681
rect -2001 647 -1985 681
rect -1885 647 -1869 681
rect -1743 647 -1727 681
rect -1627 647 -1611 681
rect -1485 647 -1469 681
rect -1369 647 -1353 681
rect -1227 647 -1211 681
rect -1111 647 -1095 681
rect -969 647 -953 681
rect -853 647 -837 681
rect -711 647 -695 681
rect -595 647 -579 681
rect -453 647 -437 681
rect -337 647 -321 681
rect -195 647 -179 681
rect -79 647 -63 681
rect 63 647 79 681
rect 179 647 195 681
rect 321 647 337 681
rect 437 647 453 681
rect 579 647 595 681
rect 695 647 711 681
rect 837 647 853 681
rect 953 647 969 681
rect 1095 647 1111 681
rect 1211 647 1227 681
rect 1353 647 1369 681
rect 1469 647 1485 681
rect 1611 647 1627 681
rect 1727 647 1743 681
rect 1869 647 1885 681
rect 1985 647 2001 681
rect 2127 647 2143 681
rect 2243 647 2259 681
rect 2385 647 2401 681
rect 2501 647 2517 681
rect 2643 647 2659 681
rect 2759 647 2775 681
rect 2901 647 2917 681
rect 3017 647 3033 681
rect 3159 647 3175 681
rect 3275 647 3291 681
rect -3371 588 -3337 604
rect -3371 -604 -3337 -588
rect -3113 588 -3079 604
rect -3113 -604 -3079 -588
rect -2855 588 -2821 604
rect -2855 -604 -2821 -588
rect -2597 588 -2563 604
rect -2597 -604 -2563 -588
rect -2339 588 -2305 604
rect -2339 -604 -2305 -588
rect -2081 588 -2047 604
rect -2081 -604 -2047 -588
rect -1823 588 -1789 604
rect -1823 -604 -1789 -588
rect -1565 588 -1531 604
rect -1565 -604 -1531 -588
rect -1307 588 -1273 604
rect -1307 -604 -1273 -588
rect -1049 588 -1015 604
rect -1049 -604 -1015 -588
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -533 588 -499 604
rect -533 -604 -499 -588
rect -275 588 -241 604
rect -275 -604 -241 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 241 588 275 604
rect 241 -604 275 -588
rect 499 588 533 604
rect 499 -604 533 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect 1015 588 1049 604
rect 1015 -604 1049 -588
rect 1273 588 1307 604
rect 1273 -604 1307 -588
rect 1531 588 1565 604
rect 1531 -604 1565 -588
rect 1789 588 1823 604
rect 1789 -604 1823 -588
rect 2047 588 2081 604
rect 2047 -604 2081 -588
rect 2305 588 2339 604
rect 2305 -604 2339 -588
rect 2563 588 2597 604
rect 2563 -604 2597 -588
rect 2821 588 2855 604
rect 2821 -604 2855 -588
rect 3079 588 3113 604
rect 3079 -604 3113 -588
rect 3337 588 3371 604
rect 3337 -604 3371 -588
rect -3291 -681 -3275 -647
rect -3175 -681 -3159 -647
rect -3033 -681 -3017 -647
rect -2917 -681 -2901 -647
rect -2775 -681 -2759 -647
rect -2659 -681 -2643 -647
rect -2517 -681 -2501 -647
rect -2401 -681 -2385 -647
rect -2259 -681 -2243 -647
rect -2143 -681 -2127 -647
rect -2001 -681 -1985 -647
rect -1885 -681 -1869 -647
rect -1743 -681 -1727 -647
rect -1627 -681 -1611 -647
rect -1485 -681 -1469 -647
rect -1369 -681 -1353 -647
rect -1227 -681 -1211 -647
rect -1111 -681 -1095 -647
rect -969 -681 -953 -647
rect -853 -681 -837 -647
rect -711 -681 -695 -647
rect -595 -681 -579 -647
rect -453 -681 -437 -647
rect -337 -681 -321 -647
rect -195 -681 -179 -647
rect -79 -681 -63 -647
rect 63 -681 79 -647
rect 179 -681 195 -647
rect 321 -681 337 -647
rect 437 -681 453 -647
rect 579 -681 595 -647
rect 695 -681 711 -647
rect 837 -681 853 -647
rect 953 -681 969 -647
rect 1095 -681 1111 -647
rect 1211 -681 1227 -647
rect 1353 -681 1369 -647
rect 1469 -681 1485 -647
rect 1611 -681 1627 -647
rect 1727 -681 1743 -647
rect 1869 -681 1885 -647
rect 1985 -681 2001 -647
rect 2127 -681 2143 -647
rect 2243 -681 2259 -647
rect 2385 -681 2401 -647
rect 2501 -681 2517 -647
rect 2643 -681 2659 -647
rect 2759 -681 2775 -647
rect 2901 -681 2917 -647
rect 3017 -681 3033 -647
rect 3159 -681 3175 -647
rect 3275 -681 3291 -647
rect -3505 -785 -3471 -723
rect 3471 -785 3505 -723
rect -3505 -819 -3409 -785
rect 3409 -819 3505 -785
<< viali >>
rect -3275 647 -3175 681
rect -3017 647 -2917 681
rect -2759 647 -2659 681
rect -2501 647 -2401 681
rect -2243 647 -2143 681
rect -1985 647 -1885 681
rect -1727 647 -1627 681
rect -1469 647 -1369 681
rect -1211 647 -1111 681
rect -953 647 -853 681
rect -695 647 -595 681
rect -437 647 -337 681
rect -179 647 -79 681
rect 79 647 179 681
rect 337 647 437 681
rect 595 647 695 681
rect 853 647 953 681
rect 1111 647 1211 681
rect 1369 647 1469 681
rect 1627 647 1727 681
rect 1885 647 1985 681
rect 2143 647 2243 681
rect 2401 647 2501 681
rect 2659 647 2759 681
rect 2917 647 3017 681
rect 3175 647 3275 681
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
rect -3275 -681 -3175 -647
rect -3017 -681 -2917 -647
rect -2759 -681 -2659 -647
rect -2501 -681 -2401 -647
rect -2243 -681 -2143 -647
rect -1985 -681 -1885 -647
rect -1727 -681 -1627 -647
rect -1469 -681 -1369 -647
rect -1211 -681 -1111 -647
rect -953 -681 -853 -647
rect -695 -681 -595 -647
rect -437 -681 -337 -647
rect -179 -681 -79 -647
rect 79 -681 179 -647
rect 337 -681 437 -647
rect 595 -681 695 -647
rect 853 -681 953 -647
rect 1111 -681 1211 -647
rect 1369 -681 1469 -647
rect 1627 -681 1727 -647
rect 1885 -681 1985 -647
rect 2143 -681 2243 -647
rect 2401 -681 2501 -647
rect 2659 -681 2759 -647
rect 2917 -681 3017 -647
rect 3175 -681 3275 -647
<< metal1 >>
rect -3287 681 -3163 687
rect -3287 647 -3275 681
rect -3175 647 -3163 681
rect -3287 641 -3163 647
rect -3029 681 -2905 687
rect -3029 647 -3017 681
rect -2917 647 -2905 681
rect -3029 641 -2905 647
rect -2771 681 -2647 687
rect -2771 647 -2759 681
rect -2659 647 -2647 681
rect -2771 641 -2647 647
rect -2513 681 -2389 687
rect -2513 647 -2501 681
rect -2401 647 -2389 681
rect -2513 641 -2389 647
rect -2255 681 -2131 687
rect -2255 647 -2243 681
rect -2143 647 -2131 681
rect -2255 641 -2131 647
rect -1997 681 -1873 687
rect -1997 647 -1985 681
rect -1885 647 -1873 681
rect -1997 641 -1873 647
rect -1739 681 -1615 687
rect -1739 647 -1727 681
rect -1627 647 -1615 681
rect -1739 641 -1615 647
rect -1481 681 -1357 687
rect -1481 647 -1469 681
rect -1369 647 -1357 681
rect -1481 641 -1357 647
rect -1223 681 -1099 687
rect -1223 647 -1211 681
rect -1111 647 -1099 681
rect -1223 641 -1099 647
rect -965 681 -841 687
rect -965 647 -953 681
rect -853 647 -841 681
rect -965 641 -841 647
rect -707 681 -583 687
rect -707 647 -695 681
rect -595 647 -583 681
rect -707 641 -583 647
rect -449 681 -325 687
rect -449 647 -437 681
rect -337 647 -325 681
rect -449 641 -325 647
rect -191 681 -67 687
rect -191 647 -179 681
rect -79 647 -67 681
rect -191 641 -67 647
rect 67 681 191 687
rect 67 647 79 681
rect 179 647 191 681
rect 67 641 191 647
rect 325 681 449 687
rect 325 647 337 681
rect 437 647 449 681
rect 325 641 449 647
rect 583 681 707 687
rect 583 647 595 681
rect 695 647 707 681
rect 583 641 707 647
rect 841 681 965 687
rect 841 647 853 681
rect 953 647 965 681
rect 841 641 965 647
rect 1099 681 1223 687
rect 1099 647 1111 681
rect 1211 647 1223 681
rect 1099 641 1223 647
rect 1357 681 1481 687
rect 1357 647 1369 681
rect 1469 647 1481 681
rect 1357 641 1481 647
rect 1615 681 1739 687
rect 1615 647 1627 681
rect 1727 647 1739 681
rect 1615 641 1739 647
rect 1873 681 1997 687
rect 1873 647 1885 681
rect 1985 647 1997 681
rect 1873 641 1997 647
rect 2131 681 2255 687
rect 2131 647 2143 681
rect 2243 647 2255 681
rect 2131 641 2255 647
rect 2389 681 2513 687
rect 2389 647 2401 681
rect 2501 647 2513 681
rect 2389 641 2513 647
rect 2647 681 2771 687
rect 2647 647 2659 681
rect 2759 647 2771 681
rect 2647 641 2771 647
rect 2905 681 3029 687
rect 2905 647 2917 681
rect 3017 647 3029 681
rect 2905 641 3029 647
rect 3163 681 3287 687
rect 3163 647 3175 681
rect 3275 647 3287 681
rect 3163 641 3287 647
rect -3377 588 -3331 600
rect -3377 -588 -3371 588
rect -3337 -588 -3331 588
rect -3377 -600 -3331 -588
rect -3119 588 -3073 600
rect -3119 -588 -3113 588
rect -3079 -588 -3073 588
rect -3119 -600 -3073 -588
rect -2861 588 -2815 600
rect -2861 -588 -2855 588
rect -2821 -588 -2815 588
rect -2861 -600 -2815 -588
rect -2603 588 -2557 600
rect -2603 -588 -2597 588
rect -2563 -588 -2557 588
rect -2603 -600 -2557 -588
rect -2345 588 -2299 600
rect -2345 -588 -2339 588
rect -2305 -588 -2299 588
rect -2345 -600 -2299 -588
rect -2087 588 -2041 600
rect -2087 -588 -2081 588
rect -2047 -588 -2041 588
rect -2087 -600 -2041 -588
rect -1829 588 -1783 600
rect -1829 -588 -1823 588
rect -1789 -588 -1783 588
rect -1829 -600 -1783 -588
rect -1571 588 -1525 600
rect -1571 -588 -1565 588
rect -1531 -588 -1525 588
rect -1571 -600 -1525 -588
rect -1313 588 -1267 600
rect -1313 -588 -1307 588
rect -1273 -588 -1267 588
rect -1313 -600 -1267 -588
rect -1055 588 -1009 600
rect -1055 -588 -1049 588
rect -1015 -588 -1009 588
rect -1055 -600 -1009 -588
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -539 588 -493 600
rect -539 -588 -533 588
rect -499 -588 -493 588
rect -539 -600 -493 -588
rect -281 588 -235 600
rect -281 -588 -275 588
rect -241 -588 -235 588
rect -281 -600 -235 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 235 588 281 600
rect 235 -588 241 588
rect 275 -588 281 588
rect 235 -600 281 -588
rect 493 588 539 600
rect 493 -588 499 588
rect 533 -588 539 588
rect 493 -600 539 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect 1009 588 1055 600
rect 1009 -588 1015 588
rect 1049 -588 1055 588
rect 1009 -600 1055 -588
rect 1267 588 1313 600
rect 1267 -588 1273 588
rect 1307 -588 1313 588
rect 1267 -600 1313 -588
rect 1525 588 1571 600
rect 1525 -588 1531 588
rect 1565 -588 1571 588
rect 1525 -600 1571 -588
rect 1783 588 1829 600
rect 1783 -588 1789 588
rect 1823 -588 1829 588
rect 1783 -600 1829 -588
rect 2041 588 2087 600
rect 2041 -588 2047 588
rect 2081 -588 2087 588
rect 2041 -600 2087 -588
rect 2299 588 2345 600
rect 2299 -588 2305 588
rect 2339 -588 2345 588
rect 2299 -600 2345 -588
rect 2557 588 2603 600
rect 2557 -588 2563 588
rect 2597 -588 2603 588
rect 2557 -600 2603 -588
rect 2815 588 2861 600
rect 2815 -588 2821 588
rect 2855 -588 2861 588
rect 2815 -600 2861 -588
rect 3073 588 3119 600
rect 3073 -588 3079 588
rect 3113 -588 3119 588
rect 3073 -600 3119 -588
rect 3331 588 3377 600
rect 3331 -588 3337 588
rect 3371 -588 3377 588
rect 3331 -600 3377 -588
rect -3287 -647 -3163 -641
rect -3287 -681 -3275 -647
rect -3175 -681 -3163 -647
rect -3287 -687 -3163 -681
rect -3029 -647 -2905 -641
rect -3029 -681 -3017 -647
rect -2917 -681 -2905 -647
rect -3029 -687 -2905 -681
rect -2771 -647 -2647 -641
rect -2771 -681 -2759 -647
rect -2659 -681 -2647 -647
rect -2771 -687 -2647 -681
rect -2513 -647 -2389 -641
rect -2513 -681 -2501 -647
rect -2401 -681 -2389 -647
rect -2513 -687 -2389 -681
rect -2255 -647 -2131 -641
rect -2255 -681 -2243 -647
rect -2143 -681 -2131 -647
rect -2255 -687 -2131 -681
rect -1997 -647 -1873 -641
rect -1997 -681 -1985 -647
rect -1885 -681 -1873 -647
rect -1997 -687 -1873 -681
rect -1739 -647 -1615 -641
rect -1739 -681 -1727 -647
rect -1627 -681 -1615 -647
rect -1739 -687 -1615 -681
rect -1481 -647 -1357 -641
rect -1481 -681 -1469 -647
rect -1369 -681 -1357 -647
rect -1481 -687 -1357 -681
rect -1223 -647 -1099 -641
rect -1223 -681 -1211 -647
rect -1111 -681 -1099 -647
rect -1223 -687 -1099 -681
rect -965 -647 -841 -641
rect -965 -681 -953 -647
rect -853 -681 -841 -647
rect -965 -687 -841 -681
rect -707 -647 -583 -641
rect -707 -681 -695 -647
rect -595 -681 -583 -647
rect -707 -687 -583 -681
rect -449 -647 -325 -641
rect -449 -681 -437 -647
rect -337 -681 -325 -647
rect -449 -687 -325 -681
rect -191 -647 -67 -641
rect -191 -681 -179 -647
rect -79 -681 -67 -647
rect -191 -687 -67 -681
rect 67 -647 191 -641
rect 67 -681 79 -647
rect 179 -681 191 -647
rect 67 -687 191 -681
rect 325 -647 449 -641
rect 325 -681 337 -647
rect 437 -681 449 -647
rect 325 -687 449 -681
rect 583 -647 707 -641
rect 583 -681 595 -647
rect 695 -681 707 -647
rect 583 -687 707 -681
rect 841 -647 965 -641
rect 841 -681 853 -647
rect 953 -681 965 -647
rect 841 -687 965 -681
rect 1099 -647 1223 -641
rect 1099 -681 1111 -647
rect 1211 -681 1223 -647
rect 1099 -687 1223 -681
rect 1357 -647 1481 -641
rect 1357 -681 1369 -647
rect 1469 -681 1481 -647
rect 1357 -687 1481 -681
rect 1615 -647 1739 -641
rect 1615 -681 1627 -647
rect 1727 -681 1739 -647
rect 1615 -687 1739 -681
rect 1873 -647 1997 -641
rect 1873 -681 1885 -647
rect 1985 -681 1997 -647
rect 1873 -687 1997 -681
rect 2131 -647 2255 -641
rect 2131 -681 2143 -647
rect 2243 -681 2255 -647
rect 2131 -687 2255 -681
rect 2389 -647 2513 -641
rect 2389 -681 2401 -647
rect 2501 -681 2513 -647
rect 2389 -687 2513 -681
rect 2647 -647 2771 -641
rect 2647 -681 2659 -647
rect 2759 -681 2771 -647
rect 2647 -687 2771 -681
rect 2905 -647 3029 -641
rect 2905 -681 2917 -647
rect 3017 -681 3029 -647
rect 2905 -687 3029 -681
rect 3163 -647 3287 -641
rect 3163 -681 3175 -647
rect 3275 -681 3287 -647
rect 3163 -687 3287 -681
<< properties >>
string FIXED_BBOX -3488 -802 3488 802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6 l 1 m 1 nf 26 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713660561
<< pwell >>
rect -584 -685 584 685
<< mvndiff >>
rect -402 491 -318 503
rect -402 457 -390 491
rect -330 457 -318 491
rect -402 400 -318 457
rect -402 -457 -318 -400
rect -402 -491 -390 -457
rect -330 -491 -318 -457
rect -402 -503 -318 -491
rect -258 491 -174 503
rect -258 457 -246 491
rect -186 457 -174 491
rect -258 400 -174 457
rect -258 -457 -174 -400
rect -258 -491 -246 -457
rect -186 -491 -174 -457
rect -258 -503 -174 -491
rect -114 491 -30 503
rect -114 457 -102 491
rect -42 457 -30 491
rect -114 400 -30 457
rect -114 -457 -30 -400
rect -114 -491 -102 -457
rect -42 -491 -30 -457
rect -114 -503 -30 -491
rect 30 491 114 503
rect 30 457 42 491
rect 102 457 114 491
rect 30 400 114 457
rect 30 -457 114 -400
rect 30 -491 42 -457
rect 102 -491 114 -457
rect 30 -503 114 -491
rect 174 491 258 503
rect 174 457 186 491
rect 246 457 258 491
rect 174 400 258 457
rect 174 -457 258 -400
rect 174 -491 186 -457
rect 246 -491 258 -457
rect 174 -503 258 -491
rect 318 491 402 503
rect 318 457 330 491
rect 390 457 402 491
rect 318 400 402 457
rect 318 -457 402 -400
rect 318 -491 330 -457
rect 390 -491 402 -457
rect 318 -503 402 -491
<< mvndiffc >>
rect -390 457 -330 491
rect -390 -491 -330 -457
rect -246 457 -186 491
rect -246 -491 -186 -457
rect -102 457 -42 491
rect -102 -491 -42 -457
rect 42 457 102 491
rect 42 -491 102 -457
rect 186 457 246 491
rect 186 -491 246 -457
rect 330 457 390 491
rect 330 -491 390 -457
<< mvpsubdiff >>
rect -548 637 548 649
rect -548 603 -440 637
rect 440 603 548 637
rect -548 591 548 603
rect -548 541 -490 591
rect -548 -541 -536 541
rect -502 -541 -490 541
rect 490 541 548 591
rect -548 -591 -490 -541
rect 490 -541 502 541
rect 536 -541 548 541
rect 490 -591 548 -541
rect -548 -603 548 -591
rect -548 -637 -440 -603
rect 440 -637 548 -603
rect -548 -649 548 -637
<< mvpsubdiffcont >>
rect -440 603 440 637
rect -536 -541 -502 541
rect 502 -541 536 541
rect -440 -637 440 -603
<< mvndiffres >>
rect -402 -400 -318 400
rect -258 -400 -174 400
rect -114 -400 -30 400
rect 30 -400 114 400
rect 174 -400 258 400
rect 318 -400 402 400
<< locali >>
rect -536 603 -440 637
rect 440 603 536 637
rect -536 541 -502 603
rect 502 541 536 603
rect -406 457 -390 491
rect -330 457 -314 491
rect -262 457 -246 491
rect -186 457 -170 491
rect -118 457 -102 491
rect -42 457 -26 491
rect 26 457 42 491
rect 102 457 118 491
rect 170 457 186 491
rect 246 457 262 491
rect 314 457 330 491
rect 390 457 406 491
rect -406 -491 -390 -457
rect -330 -491 -314 -457
rect -262 -491 -246 -457
rect -186 -491 -170 -457
rect -118 -491 -102 -457
rect -42 -491 -26 -457
rect 26 -491 42 -457
rect 102 -491 118 -457
rect 170 -491 186 -457
rect 246 -491 262 -457
rect 314 -491 330 -457
rect 390 -491 406 -457
rect -536 -603 -502 -541
rect 502 -603 536 -541
rect -536 -637 -440 -603
rect 440 -637 536 -603
<< viali >>
rect -390 457 -330 491
rect -246 457 -186 491
rect -102 457 -42 491
rect 42 457 102 491
rect 186 457 246 491
rect 330 457 390 491
rect -390 417 -330 457
rect -246 417 -186 457
rect -102 417 -42 457
rect 42 417 102 457
rect 186 417 246 457
rect 330 417 390 457
rect -390 -457 -330 -417
rect -246 -457 -186 -417
rect -102 -457 -42 -417
rect 42 -457 102 -417
rect 186 -457 246 -417
rect 330 -457 390 -417
rect -390 -491 -330 -457
rect -246 -491 -186 -457
rect -102 -491 -42 -457
rect 42 -491 102 -457
rect 186 -491 246 -457
rect 330 -491 390 -457
<< metal1 >>
rect -396 491 -324 503
rect -396 417 -390 491
rect -330 417 -324 491
rect -396 405 -324 417
rect -252 491 -180 503
rect -252 417 -246 491
rect -186 417 -180 491
rect -252 405 -180 417
rect -108 491 -36 503
rect -108 417 -102 491
rect -42 417 -36 491
rect -108 405 -36 417
rect 36 491 108 503
rect 36 417 42 491
rect 102 417 108 491
rect 36 405 108 417
rect 180 491 252 503
rect 180 417 186 491
rect 246 417 252 491
rect 180 405 252 417
rect 324 491 396 503
rect 324 417 330 491
rect 390 417 396 491
rect 324 405 396 417
rect -396 -417 -324 -405
rect -396 -491 -390 -417
rect -330 -491 -324 -417
rect -396 -503 -324 -491
rect -252 -417 -180 -405
rect -252 -491 -246 -417
rect -186 -491 -180 -417
rect -252 -503 -180 -491
rect -108 -417 -36 -405
rect -108 -491 -102 -417
rect -42 -491 -36 -417
rect -108 -503 -36 -491
rect 36 -417 108 -405
rect 36 -491 42 -417
rect 102 -491 108 -417
rect 36 -503 108 -491
rect 180 -417 252 -405
rect 180 -491 186 -417
rect 246 -491 252 -417
rect 180 -503 252 -491
rect 324 -417 396 -405
rect 324 -491 330 -417
rect 390 -491 396 -417
rect 324 -503 396 -491
<< properties >>
string FIXED_BBOX -519 -620 519 620
string gencell sky130_fd_pr__res_generic_nd__hv
string library sky130
string parameters w 0.420 l 4 m 1 nx 6 wmin 0.42 lmin 2.10 rho 120 val 1.2k dummy 0 dw 0.02 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713300479
<< error_p >>
rect -743 522 -679 528
rect -585 522 -521 528
rect -427 522 -363 528
rect -269 522 -205 528
rect -111 522 -47 528
rect 47 522 111 528
rect 205 522 269 528
rect 363 522 427 528
rect 521 522 585 528
rect 679 522 743 528
rect -743 488 -731 522
rect -585 488 -573 522
rect -427 488 -415 522
rect -269 488 -257 522
rect -111 488 -99 522
rect 47 488 59 522
rect 205 488 217 522
rect 363 488 375 522
rect 521 488 533 522
rect 679 488 691 522
rect -743 482 -679 488
rect -585 482 -521 488
rect -427 482 -363 488
rect -269 482 -205 488
rect -111 482 -47 488
rect 47 482 111 488
rect 205 482 269 488
rect 363 482 427 488
rect 521 482 585 488
rect 679 482 743 488
rect -743 -488 -679 -482
rect -585 -488 -521 -482
rect -427 -488 -363 -482
rect -269 -488 -205 -482
rect -111 -488 -47 -482
rect 47 -488 111 -482
rect 205 -488 269 -482
rect 363 -488 427 -482
rect 521 -488 585 -482
rect 679 -488 743 -482
rect -743 -522 -731 -488
rect -585 -522 -573 -488
rect -427 -522 -415 -488
rect -269 -522 -257 -488
rect -111 -522 -99 -488
rect 47 -522 59 -488
rect 205 -522 217 -488
rect 363 -522 375 -488
rect 521 -522 533 -488
rect 679 -522 691 -488
rect -743 -528 -679 -522
rect -585 -528 -521 -522
rect -427 -528 -363 -522
rect -269 -528 -205 -522
rect -111 -528 -47 -522
rect 47 -528 111 -522
rect 205 -528 269 -522
rect 363 -528 427 -522
rect 521 -528 585 -522
rect 679 -528 743 -522
<< pwell >>
rect -989 -708 989 708
<< mvnmos >>
rect -761 -450 -661 450
rect -603 -450 -503 450
rect -445 -450 -345 450
rect -287 -450 -187 450
rect -129 -450 -29 450
rect 29 -450 129 450
rect 187 -450 287 450
rect 345 -450 445 450
rect 503 -450 603 450
rect 661 -450 761 450
<< mvndiff >>
rect -819 438 -761 450
rect -819 -438 -807 438
rect -773 -438 -761 438
rect -819 -450 -761 -438
rect -661 438 -603 450
rect -661 -438 -649 438
rect -615 -438 -603 438
rect -661 -450 -603 -438
rect -503 438 -445 450
rect -503 -438 -491 438
rect -457 -438 -445 438
rect -503 -450 -445 -438
rect -345 438 -287 450
rect -345 -438 -333 438
rect -299 -438 -287 438
rect -345 -450 -287 -438
rect -187 438 -129 450
rect -187 -438 -175 438
rect -141 -438 -129 438
rect -187 -450 -129 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 129 438 187 450
rect 129 -438 141 438
rect 175 -438 187 438
rect 129 -450 187 -438
rect 287 438 345 450
rect 287 -438 299 438
rect 333 -438 345 438
rect 287 -450 345 -438
rect 445 438 503 450
rect 445 -438 457 438
rect 491 -438 503 438
rect 445 -450 503 -438
rect 603 438 661 450
rect 603 -438 615 438
rect 649 -438 661 438
rect 603 -450 661 -438
rect 761 438 819 450
rect 761 -438 773 438
rect 807 -438 819 438
rect 761 -450 819 -438
<< mvndiffc >>
rect -807 -438 -773 438
rect -649 -438 -615 438
rect -491 -438 -457 438
rect -333 -438 -299 438
rect -175 -438 -141 438
rect -17 -438 17 438
rect 141 -438 175 438
rect 299 -438 333 438
rect 457 -438 491 438
rect 615 -438 649 438
rect 773 -438 807 438
<< mvpsubdiff >>
rect -953 660 953 672
rect -953 626 -845 660
rect 845 626 953 660
rect -953 614 953 626
rect -953 564 -895 614
rect -953 -564 -941 564
rect -907 -564 -895 564
rect 895 564 953 614
rect -953 -614 -895 -564
rect 895 -564 907 564
rect 941 -564 953 564
rect 895 -614 953 -564
rect -953 -626 953 -614
rect -953 -660 -845 -626
rect 845 -660 953 -626
rect -953 -672 953 -660
<< mvpsubdiffcont >>
rect -845 626 845 660
rect -941 -564 -907 564
rect 907 -564 941 564
rect -845 -660 845 -626
<< poly >>
rect -747 522 -675 538
rect -747 505 -731 522
rect -761 488 -731 505
rect -691 505 -675 522
rect -589 522 -517 538
rect -589 505 -573 522
rect -691 488 -661 505
rect -761 450 -661 488
rect -603 488 -573 505
rect -533 505 -517 522
rect -431 522 -359 538
rect -431 505 -415 522
rect -533 488 -503 505
rect -603 450 -503 488
rect -445 488 -415 505
rect -375 505 -359 522
rect -273 522 -201 538
rect -273 505 -257 522
rect -375 488 -345 505
rect -445 450 -345 488
rect -287 488 -257 505
rect -217 505 -201 522
rect -115 522 -43 538
rect -115 505 -99 522
rect -217 488 -187 505
rect -287 450 -187 488
rect -129 488 -99 505
rect -59 505 -43 522
rect 43 522 115 538
rect 43 505 59 522
rect -59 488 -29 505
rect -129 450 -29 488
rect 29 488 59 505
rect 99 505 115 522
rect 201 522 273 538
rect 201 505 217 522
rect 99 488 129 505
rect 29 450 129 488
rect 187 488 217 505
rect 257 505 273 522
rect 359 522 431 538
rect 359 505 375 522
rect 257 488 287 505
rect 187 450 287 488
rect 345 488 375 505
rect 415 505 431 522
rect 517 522 589 538
rect 517 505 533 522
rect 415 488 445 505
rect 345 450 445 488
rect 503 488 533 505
rect 573 505 589 522
rect 675 522 747 538
rect 675 505 691 522
rect 573 488 603 505
rect 503 450 603 488
rect 661 488 691 505
rect 731 505 747 522
rect 731 488 761 505
rect 661 450 761 488
rect -761 -488 -661 -450
rect -761 -505 -731 -488
rect -747 -522 -731 -505
rect -691 -505 -661 -488
rect -603 -488 -503 -450
rect -603 -505 -573 -488
rect -691 -522 -675 -505
rect -747 -538 -675 -522
rect -589 -522 -573 -505
rect -533 -505 -503 -488
rect -445 -488 -345 -450
rect -445 -505 -415 -488
rect -533 -522 -517 -505
rect -589 -538 -517 -522
rect -431 -522 -415 -505
rect -375 -505 -345 -488
rect -287 -488 -187 -450
rect -287 -505 -257 -488
rect -375 -522 -359 -505
rect -431 -538 -359 -522
rect -273 -522 -257 -505
rect -217 -505 -187 -488
rect -129 -488 -29 -450
rect -129 -505 -99 -488
rect -217 -522 -201 -505
rect -273 -538 -201 -522
rect -115 -522 -99 -505
rect -59 -505 -29 -488
rect 29 -488 129 -450
rect 29 -505 59 -488
rect -59 -522 -43 -505
rect -115 -538 -43 -522
rect 43 -522 59 -505
rect 99 -505 129 -488
rect 187 -488 287 -450
rect 187 -505 217 -488
rect 99 -522 115 -505
rect 43 -538 115 -522
rect 201 -522 217 -505
rect 257 -505 287 -488
rect 345 -488 445 -450
rect 345 -505 375 -488
rect 257 -522 273 -505
rect 201 -538 273 -522
rect 359 -522 375 -505
rect 415 -505 445 -488
rect 503 -488 603 -450
rect 503 -505 533 -488
rect 415 -522 431 -505
rect 359 -538 431 -522
rect 517 -522 533 -505
rect 573 -505 603 -488
rect 661 -488 761 -450
rect 661 -505 691 -488
rect 573 -522 589 -505
rect 517 -538 589 -522
rect 675 -522 691 -505
rect 731 -505 761 -488
rect 731 -522 747 -505
rect 675 -538 747 -522
<< polycont >>
rect -731 488 -691 522
rect -573 488 -533 522
rect -415 488 -375 522
rect -257 488 -217 522
rect -99 488 -59 522
rect 59 488 99 522
rect 217 488 257 522
rect 375 488 415 522
rect 533 488 573 522
rect 691 488 731 522
rect -731 -522 -691 -488
rect -573 -522 -533 -488
rect -415 -522 -375 -488
rect -257 -522 -217 -488
rect -99 -522 -59 -488
rect 59 -522 99 -488
rect 217 -522 257 -488
rect 375 -522 415 -488
rect 533 -522 573 -488
rect 691 -522 731 -488
<< locali >>
rect -941 626 -845 660
rect 845 626 941 660
rect -941 564 -907 626
rect 907 564 941 626
rect -747 488 -731 522
rect -691 488 -675 522
rect -589 488 -573 522
rect -533 488 -517 522
rect -431 488 -415 522
rect -375 488 -359 522
rect -273 488 -257 522
rect -217 488 -201 522
rect -115 488 -99 522
rect -59 488 -43 522
rect 43 488 59 522
rect 99 488 115 522
rect 201 488 217 522
rect 257 488 273 522
rect 359 488 375 522
rect 415 488 431 522
rect 517 488 533 522
rect 573 488 589 522
rect 675 488 691 522
rect 731 488 747 522
rect -807 438 -773 454
rect -807 -454 -773 -438
rect -649 438 -615 454
rect -649 -454 -615 -438
rect -491 438 -457 454
rect -491 -454 -457 -438
rect -333 438 -299 454
rect -333 -454 -299 -438
rect -175 438 -141 454
rect -175 -454 -141 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 141 438 175 454
rect 141 -454 175 -438
rect 299 438 333 454
rect 299 -454 333 -438
rect 457 438 491 454
rect 457 -454 491 -438
rect 615 438 649 454
rect 615 -454 649 -438
rect 773 438 807 454
rect 773 -454 807 -438
rect -747 -522 -731 -488
rect -691 -522 -675 -488
rect -589 -522 -573 -488
rect -533 -522 -517 -488
rect -431 -522 -415 -488
rect -375 -522 -359 -488
rect -273 -522 -257 -488
rect -217 -522 -201 -488
rect -115 -522 -99 -488
rect -59 -522 -43 -488
rect 43 -522 59 -488
rect 99 -522 115 -488
rect 201 -522 217 -488
rect 257 -522 273 -488
rect 359 -522 375 -488
rect 415 -522 431 -488
rect 517 -522 533 -488
rect 573 -522 589 -488
rect 675 -522 691 -488
rect 731 -522 747 -488
rect -941 -626 -907 -564
rect 907 -626 941 -564
rect -941 -660 -845 -626
rect 845 -660 941 -626
<< viali >>
rect -731 488 -691 522
rect -573 488 -533 522
rect -415 488 -375 522
rect -257 488 -217 522
rect -99 488 -59 522
rect 59 488 99 522
rect 217 488 257 522
rect 375 488 415 522
rect 533 488 573 522
rect 691 488 731 522
rect -807 -438 -773 438
rect -649 -438 -615 438
rect -491 -438 -457 438
rect -333 -438 -299 438
rect -175 -438 -141 438
rect -17 -438 17 438
rect 141 -438 175 438
rect 299 -438 333 438
rect 457 -438 491 438
rect 615 -438 649 438
rect 773 -438 807 438
rect -731 -522 -691 -488
rect -573 -522 -533 -488
rect -415 -522 -375 -488
rect -257 -522 -217 -488
rect -99 -522 -59 -488
rect 59 -522 99 -488
rect 217 -522 257 -488
rect 375 -522 415 -488
rect 533 -522 573 -488
rect 691 -522 731 -488
<< metal1 >>
rect -743 522 -679 528
rect -743 488 -731 522
rect -691 488 -679 522
rect -743 482 -679 488
rect -585 522 -521 528
rect -585 488 -573 522
rect -533 488 -521 522
rect -585 482 -521 488
rect -427 522 -363 528
rect -427 488 -415 522
rect -375 488 -363 522
rect -427 482 -363 488
rect -269 522 -205 528
rect -269 488 -257 522
rect -217 488 -205 522
rect -269 482 -205 488
rect -111 522 -47 528
rect -111 488 -99 522
rect -59 488 -47 522
rect -111 482 -47 488
rect 47 522 111 528
rect 47 488 59 522
rect 99 488 111 522
rect 47 482 111 488
rect 205 522 269 528
rect 205 488 217 522
rect 257 488 269 522
rect 205 482 269 488
rect 363 522 427 528
rect 363 488 375 522
rect 415 488 427 522
rect 363 482 427 488
rect 521 522 585 528
rect 521 488 533 522
rect 573 488 585 522
rect 521 482 585 488
rect 679 522 743 528
rect 679 488 691 522
rect 731 488 743 522
rect 679 482 743 488
rect -813 438 -767 450
rect -813 -438 -807 438
rect -773 -438 -767 438
rect -813 -450 -767 -438
rect -655 438 -609 450
rect -655 -438 -649 438
rect -615 -438 -609 438
rect -655 -450 -609 -438
rect -497 438 -451 450
rect -497 -438 -491 438
rect -457 -438 -451 438
rect -497 -450 -451 -438
rect -339 438 -293 450
rect -339 -438 -333 438
rect -299 -438 -293 438
rect -339 -450 -293 -438
rect -181 438 -135 450
rect -181 -438 -175 438
rect -141 -438 -135 438
rect -181 -450 -135 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 135 438 181 450
rect 135 -438 141 438
rect 175 -438 181 438
rect 135 -450 181 -438
rect 293 438 339 450
rect 293 -438 299 438
rect 333 -438 339 438
rect 293 -450 339 -438
rect 451 438 497 450
rect 451 -438 457 438
rect 491 -438 497 438
rect 451 -450 497 -438
rect 609 438 655 450
rect 609 -438 615 438
rect 649 -438 655 438
rect 609 -450 655 -438
rect 767 438 813 450
rect 767 -438 773 438
rect 807 -438 813 438
rect 767 -450 813 -438
rect -743 -488 -679 -482
rect -743 -522 -731 -488
rect -691 -522 -679 -488
rect -743 -528 -679 -522
rect -585 -488 -521 -482
rect -585 -522 -573 -488
rect -533 -522 -521 -488
rect -585 -528 -521 -522
rect -427 -488 -363 -482
rect -427 -522 -415 -488
rect -375 -522 -363 -488
rect -427 -528 -363 -522
rect -269 -488 -205 -482
rect -269 -522 -257 -488
rect -217 -522 -205 -488
rect -269 -528 -205 -522
rect -111 -488 -47 -482
rect -111 -522 -99 -488
rect -59 -522 -47 -488
rect -111 -528 -47 -522
rect 47 -488 111 -482
rect 47 -522 59 -488
rect 99 -522 111 -488
rect 47 -528 111 -522
rect 205 -488 269 -482
rect 205 -522 217 -488
rect 257 -522 269 -488
rect 205 -528 269 -522
rect 363 -488 427 -482
rect 363 -522 375 -488
rect 415 -522 427 -488
rect 363 -528 427 -522
rect 521 -488 585 -482
rect 521 -522 533 -488
rect 573 -522 585 -488
rect 521 -528 585 -522
rect 679 -488 743 -482
rect 679 -522 691 -488
rect 731 -522 743 -488
rect 679 -528 743 -522
<< properties >>
string FIXED_BBOX -924 -643 924 643
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 0.5 m 1 nf 10 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

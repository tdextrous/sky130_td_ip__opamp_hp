magic
tech sky130A
magscale 1 2
timestamp 1713331128
<< nwell >>
rect -1777 -497 1777 497
<< mvpmos >>
rect -1519 -200 -1319 200
rect -1261 -200 -1061 200
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
rect 1061 -200 1261 200
rect 1319 -200 1519 200
<< mvpdiff >>
rect -1577 188 -1519 200
rect -1577 -188 -1565 188
rect -1531 -188 -1519 188
rect -1577 -200 -1519 -188
rect -1319 188 -1261 200
rect -1319 -188 -1307 188
rect -1273 -188 -1261 188
rect -1319 -200 -1261 -188
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
rect 1261 188 1319 200
rect 1261 -188 1273 188
rect 1307 -188 1319 188
rect 1261 -200 1319 -188
rect 1519 188 1577 200
rect 1519 -188 1531 188
rect 1565 -188 1577 188
rect 1519 -200 1577 -188
<< mvpdiffc >>
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
<< mvnsubdiff >>
rect -1711 419 1711 431
rect -1711 385 -1603 419
rect 1603 385 1711 419
rect -1711 373 1711 385
rect -1711 323 -1653 373
rect -1711 -323 -1699 323
rect -1665 -323 -1653 323
rect 1653 323 1711 373
rect -1711 -373 -1653 -323
rect 1653 -323 1665 323
rect 1699 -323 1711 323
rect 1653 -373 1711 -323
rect -1711 -385 1711 -373
rect -1711 -419 -1603 -385
rect 1603 -419 1711 -385
rect -1711 -431 1711 -419
<< mvnsubdiffcont >>
rect -1603 385 1603 419
rect -1699 -323 -1665 323
rect 1665 -323 1699 323
rect -1603 -419 1603 -385
<< poly >>
rect -1485 281 -1353 297
rect -1485 264 -1469 281
rect -1519 247 -1469 264
rect -1369 264 -1353 281
rect -1227 281 -1095 297
rect -1227 264 -1211 281
rect -1369 247 -1319 264
rect -1519 200 -1319 247
rect -1261 247 -1211 264
rect -1111 264 -1095 281
rect -969 281 -837 297
rect -969 264 -953 281
rect -1111 247 -1061 264
rect -1261 200 -1061 247
rect -1003 247 -953 264
rect -853 264 -837 281
rect -711 281 -579 297
rect -711 264 -695 281
rect -853 247 -803 264
rect -1003 200 -803 247
rect -745 247 -695 264
rect -595 264 -579 281
rect -453 281 -321 297
rect -453 264 -437 281
rect -595 247 -545 264
rect -745 200 -545 247
rect -487 247 -437 264
rect -337 264 -321 281
rect -195 281 -63 297
rect -195 264 -179 281
rect -337 247 -287 264
rect -487 200 -287 247
rect -229 247 -179 264
rect -79 264 -63 281
rect 63 281 195 297
rect 63 264 79 281
rect -79 247 -29 264
rect -229 200 -29 247
rect 29 247 79 264
rect 179 264 195 281
rect 321 281 453 297
rect 321 264 337 281
rect 179 247 229 264
rect 29 200 229 247
rect 287 247 337 264
rect 437 264 453 281
rect 579 281 711 297
rect 579 264 595 281
rect 437 247 487 264
rect 287 200 487 247
rect 545 247 595 264
rect 695 264 711 281
rect 837 281 969 297
rect 837 264 853 281
rect 695 247 745 264
rect 545 200 745 247
rect 803 247 853 264
rect 953 264 969 281
rect 1095 281 1227 297
rect 1095 264 1111 281
rect 953 247 1003 264
rect 803 200 1003 247
rect 1061 247 1111 264
rect 1211 264 1227 281
rect 1353 281 1485 297
rect 1353 264 1369 281
rect 1211 247 1261 264
rect 1061 200 1261 247
rect 1319 247 1369 264
rect 1469 264 1485 281
rect 1469 247 1519 264
rect 1319 200 1519 247
rect -1519 -247 -1319 -200
rect -1519 -264 -1469 -247
rect -1485 -281 -1469 -264
rect -1369 -264 -1319 -247
rect -1261 -247 -1061 -200
rect -1261 -264 -1211 -247
rect -1369 -281 -1353 -264
rect -1485 -297 -1353 -281
rect -1227 -281 -1211 -264
rect -1111 -264 -1061 -247
rect -1003 -247 -803 -200
rect -1003 -264 -953 -247
rect -1111 -281 -1095 -264
rect -1227 -297 -1095 -281
rect -969 -281 -953 -264
rect -853 -264 -803 -247
rect -745 -247 -545 -200
rect -745 -264 -695 -247
rect -853 -281 -837 -264
rect -969 -297 -837 -281
rect -711 -281 -695 -264
rect -595 -264 -545 -247
rect -487 -247 -287 -200
rect -487 -264 -437 -247
rect -595 -281 -579 -264
rect -711 -297 -579 -281
rect -453 -281 -437 -264
rect -337 -264 -287 -247
rect -229 -247 -29 -200
rect -229 -264 -179 -247
rect -337 -281 -321 -264
rect -453 -297 -321 -281
rect -195 -281 -179 -264
rect -79 -264 -29 -247
rect 29 -247 229 -200
rect 29 -264 79 -247
rect -79 -281 -63 -264
rect -195 -297 -63 -281
rect 63 -281 79 -264
rect 179 -264 229 -247
rect 287 -247 487 -200
rect 287 -264 337 -247
rect 179 -281 195 -264
rect 63 -297 195 -281
rect 321 -281 337 -264
rect 437 -264 487 -247
rect 545 -247 745 -200
rect 545 -264 595 -247
rect 437 -281 453 -264
rect 321 -297 453 -281
rect 579 -281 595 -264
rect 695 -264 745 -247
rect 803 -247 1003 -200
rect 803 -264 853 -247
rect 695 -281 711 -264
rect 579 -297 711 -281
rect 837 -281 853 -264
rect 953 -264 1003 -247
rect 1061 -247 1261 -200
rect 1061 -264 1111 -247
rect 953 -281 969 -264
rect 837 -297 969 -281
rect 1095 -281 1111 -264
rect 1211 -264 1261 -247
rect 1319 -247 1519 -200
rect 1319 -264 1369 -247
rect 1211 -281 1227 -264
rect 1095 -297 1227 -281
rect 1353 -281 1369 -264
rect 1469 -264 1519 -247
rect 1469 -281 1485 -264
rect 1353 -297 1485 -281
<< polycont >>
rect -1469 247 -1369 281
rect -1211 247 -1111 281
rect -953 247 -853 281
rect -695 247 -595 281
rect -437 247 -337 281
rect -179 247 -79 281
rect 79 247 179 281
rect 337 247 437 281
rect 595 247 695 281
rect 853 247 953 281
rect 1111 247 1211 281
rect 1369 247 1469 281
rect -1469 -281 -1369 -247
rect -1211 -281 -1111 -247
rect -953 -281 -853 -247
rect -695 -281 -595 -247
rect -437 -281 -337 -247
rect -179 -281 -79 -247
rect 79 -281 179 -247
rect 337 -281 437 -247
rect 595 -281 695 -247
rect 853 -281 953 -247
rect 1111 -281 1211 -247
rect 1369 -281 1469 -247
<< locali >>
rect -1699 385 -1603 419
rect 1603 385 1699 419
rect -1699 323 -1665 385
rect 1665 323 1699 385
rect -1485 247 -1469 281
rect -1369 247 -1353 281
rect -1227 247 -1211 281
rect -1111 247 -1095 281
rect -969 247 -953 281
rect -853 247 -837 281
rect -711 247 -695 281
rect -595 247 -579 281
rect -453 247 -437 281
rect -337 247 -321 281
rect -195 247 -179 281
rect -79 247 -63 281
rect 63 247 79 281
rect 179 247 195 281
rect 321 247 337 281
rect 437 247 453 281
rect 579 247 595 281
rect 695 247 711 281
rect 837 247 853 281
rect 953 247 969 281
rect 1095 247 1111 281
rect 1211 247 1227 281
rect 1353 247 1369 281
rect 1469 247 1485 281
rect -1565 188 -1531 204
rect -1565 -204 -1531 -188
rect -1307 188 -1273 204
rect -1307 -204 -1273 -188
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect 1273 188 1307 204
rect 1273 -204 1307 -188
rect 1531 188 1565 204
rect 1531 -204 1565 -188
rect -1485 -281 -1469 -247
rect -1369 -281 -1353 -247
rect -1227 -281 -1211 -247
rect -1111 -281 -1095 -247
rect -969 -281 -953 -247
rect -853 -281 -837 -247
rect -711 -281 -695 -247
rect -595 -281 -579 -247
rect -453 -281 -437 -247
rect -337 -281 -321 -247
rect -195 -281 -179 -247
rect -79 -281 -63 -247
rect 63 -281 79 -247
rect 179 -281 195 -247
rect 321 -281 337 -247
rect 437 -281 453 -247
rect 579 -281 595 -247
rect 695 -281 711 -247
rect 837 -281 853 -247
rect 953 -281 969 -247
rect 1095 -281 1111 -247
rect 1211 -281 1227 -247
rect 1353 -281 1369 -247
rect 1469 -281 1485 -247
rect -1699 -385 -1665 -323
rect 1665 -385 1699 -323
rect -1699 -419 -1603 -385
rect 1603 -419 1699 -385
<< viali >>
rect -1469 247 -1369 281
rect -1211 247 -1111 281
rect -953 247 -853 281
rect -695 247 -595 281
rect -437 247 -337 281
rect -179 247 -79 281
rect 79 247 179 281
rect 337 247 437 281
rect 595 247 695 281
rect 853 247 953 281
rect 1111 247 1211 281
rect 1369 247 1469 281
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect -1469 -281 -1369 -247
rect -1211 -281 -1111 -247
rect -953 -281 -853 -247
rect -695 -281 -595 -247
rect -437 -281 -337 -247
rect -179 -281 -79 -247
rect 79 -281 179 -247
rect 337 -281 437 -247
rect 595 -281 695 -247
rect 853 -281 953 -247
rect 1111 -281 1211 -247
rect 1369 -281 1469 -247
<< metal1 >>
rect -1481 281 -1357 287
rect -1481 247 -1469 281
rect -1369 247 -1357 281
rect -1481 241 -1357 247
rect -1223 281 -1099 287
rect -1223 247 -1211 281
rect -1111 247 -1099 281
rect -1223 241 -1099 247
rect -965 281 -841 287
rect -965 247 -953 281
rect -853 247 -841 281
rect -965 241 -841 247
rect -707 281 -583 287
rect -707 247 -695 281
rect -595 247 -583 281
rect -707 241 -583 247
rect -449 281 -325 287
rect -449 247 -437 281
rect -337 247 -325 281
rect -449 241 -325 247
rect -191 281 -67 287
rect -191 247 -179 281
rect -79 247 -67 281
rect -191 241 -67 247
rect 67 281 191 287
rect 67 247 79 281
rect 179 247 191 281
rect 67 241 191 247
rect 325 281 449 287
rect 325 247 337 281
rect 437 247 449 281
rect 325 241 449 247
rect 583 281 707 287
rect 583 247 595 281
rect 695 247 707 281
rect 583 241 707 247
rect 841 281 965 287
rect 841 247 853 281
rect 953 247 965 281
rect 841 241 965 247
rect 1099 281 1223 287
rect 1099 247 1111 281
rect 1211 247 1223 281
rect 1099 241 1223 247
rect 1357 281 1481 287
rect 1357 247 1369 281
rect 1469 247 1481 281
rect 1357 241 1481 247
rect -1571 188 -1525 200
rect -1571 -188 -1565 188
rect -1531 -188 -1525 188
rect -1571 -200 -1525 -188
rect -1313 188 -1267 200
rect -1313 -188 -1307 188
rect -1273 -188 -1267 188
rect -1313 -200 -1267 -188
rect -1055 188 -1009 200
rect -1055 -188 -1049 188
rect -1015 -188 -1009 188
rect -1055 -200 -1009 -188
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect 1009 188 1055 200
rect 1009 -188 1015 188
rect 1049 -188 1055 188
rect 1009 -200 1055 -188
rect 1267 188 1313 200
rect 1267 -188 1273 188
rect 1307 -188 1313 188
rect 1267 -200 1313 -188
rect 1525 188 1571 200
rect 1525 -188 1531 188
rect 1565 -188 1571 188
rect 1525 -200 1571 -188
rect -1481 -247 -1357 -241
rect -1481 -281 -1469 -247
rect -1369 -281 -1357 -247
rect -1481 -287 -1357 -281
rect -1223 -247 -1099 -241
rect -1223 -281 -1211 -247
rect -1111 -281 -1099 -247
rect -1223 -287 -1099 -281
rect -965 -247 -841 -241
rect -965 -281 -953 -247
rect -853 -281 -841 -247
rect -965 -287 -841 -281
rect -707 -247 -583 -241
rect -707 -281 -695 -247
rect -595 -281 -583 -247
rect -707 -287 -583 -281
rect -449 -247 -325 -241
rect -449 -281 -437 -247
rect -337 -281 -325 -247
rect -449 -287 -325 -281
rect -191 -247 -67 -241
rect -191 -281 -179 -247
rect -79 -281 -67 -247
rect -191 -287 -67 -281
rect 67 -247 191 -241
rect 67 -281 79 -247
rect 179 -281 191 -247
rect 67 -287 191 -281
rect 325 -247 449 -241
rect 325 -281 337 -247
rect 437 -281 449 -247
rect 325 -287 449 -281
rect 583 -247 707 -241
rect 583 -281 595 -247
rect 695 -281 707 -247
rect 583 -287 707 -281
rect 841 -247 965 -241
rect 841 -281 853 -247
rect 953 -281 965 -247
rect 841 -287 965 -281
rect 1099 -247 1223 -241
rect 1099 -281 1111 -247
rect 1211 -281 1223 -247
rect 1099 -287 1223 -281
rect 1357 -247 1481 -241
rect 1357 -281 1369 -247
rect 1469 -281 1481 -247
rect 1357 -287 1481 -281
<< properties >>
string FIXED_BBOX -1682 -402 1682 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 12 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713393095
<< nwell >>
rect -1777 -697 1777 697
<< mvpmos >>
rect -1519 -400 -1319 400
rect -1261 -400 -1061 400
rect -1003 -400 -803 400
rect -745 -400 -545 400
rect -487 -400 -287 400
rect -229 -400 -29 400
rect 29 -400 229 400
rect 287 -400 487 400
rect 545 -400 745 400
rect 803 -400 1003 400
rect 1061 -400 1261 400
rect 1319 -400 1519 400
<< mvpdiff >>
rect -1577 388 -1519 400
rect -1577 -388 -1565 388
rect -1531 -388 -1519 388
rect -1577 -400 -1519 -388
rect -1319 388 -1261 400
rect -1319 -388 -1307 388
rect -1273 -388 -1261 388
rect -1319 -400 -1261 -388
rect -1061 388 -1003 400
rect -1061 -388 -1049 388
rect -1015 -388 -1003 388
rect -1061 -400 -1003 -388
rect -803 388 -745 400
rect -803 -388 -791 388
rect -757 -388 -745 388
rect -803 -400 -745 -388
rect -545 388 -487 400
rect -545 -388 -533 388
rect -499 -388 -487 388
rect -545 -400 -487 -388
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect 487 388 545 400
rect 487 -388 499 388
rect 533 -388 545 388
rect 487 -400 545 -388
rect 745 388 803 400
rect 745 -388 757 388
rect 791 -388 803 388
rect 745 -400 803 -388
rect 1003 388 1061 400
rect 1003 -388 1015 388
rect 1049 -388 1061 388
rect 1003 -400 1061 -388
rect 1261 388 1319 400
rect 1261 -388 1273 388
rect 1307 -388 1319 388
rect 1261 -400 1319 -388
rect 1519 388 1577 400
rect 1519 -388 1531 388
rect 1565 -388 1577 388
rect 1519 -400 1577 -388
<< mvpdiffc >>
rect -1565 -388 -1531 388
rect -1307 -388 -1273 388
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect 1273 -388 1307 388
rect 1531 -388 1565 388
<< mvnsubdiff >>
rect -1711 619 1711 631
rect -1711 585 -1603 619
rect 1603 585 1711 619
rect -1711 573 1711 585
rect -1711 523 -1653 573
rect -1711 -523 -1699 523
rect -1665 -523 -1653 523
rect 1653 523 1711 573
rect -1711 -573 -1653 -523
rect 1653 -523 1665 523
rect 1699 -523 1711 523
rect 1653 -573 1711 -523
rect -1711 -585 1711 -573
rect -1711 -619 -1603 -585
rect 1603 -619 1711 -585
rect -1711 -631 1711 -619
<< mvnsubdiffcont >>
rect -1603 585 1603 619
rect -1699 -523 -1665 523
rect 1665 -523 1699 523
rect -1603 -619 1603 -585
<< poly >>
rect -1485 481 -1353 497
rect -1485 464 -1469 481
rect -1519 447 -1469 464
rect -1369 464 -1353 481
rect -1227 481 -1095 497
rect -1227 464 -1211 481
rect -1369 447 -1319 464
rect -1519 400 -1319 447
rect -1261 447 -1211 464
rect -1111 464 -1095 481
rect -969 481 -837 497
rect -969 464 -953 481
rect -1111 447 -1061 464
rect -1261 400 -1061 447
rect -1003 447 -953 464
rect -853 464 -837 481
rect -711 481 -579 497
rect -711 464 -695 481
rect -853 447 -803 464
rect -1003 400 -803 447
rect -745 447 -695 464
rect -595 464 -579 481
rect -453 481 -321 497
rect -453 464 -437 481
rect -595 447 -545 464
rect -745 400 -545 447
rect -487 447 -437 464
rect -337 464 -321 481
rect -195 481 -63 497
rect -195 464 -179 481
rect -337 447 -287 464
rect -487 400 -287 447
rect -229 447 -179 464
rect -79 464 -63 481
rect 63 481 195 497
rect 63 464 79 481
rect -79 447 -29 464
rect -229 400 -29 447
rect 29 447 79 464
rect 179 464 195 481
rect 321 481 453 497
rect 321 464 337 481
rect 179 447 229 464
rect 29 400 229 447
rect 287 447 337 464
rect 437 464 453 481
rect 579 481 711 497
rect 579 464 595 481
rect 437 447 487 464
rect 287 400 487 447
rect 545 447 595 464
rect 695 464 711 481
rect 837 481 969 497
rect 837 464 853 481
rect 695 447 745 464
rect 545 400 745 447
rect 803 447 853 464
rect 953 464 969 481
rect 1095 481 1227 497
rect 1095 464 1111 481
rect 953 447 1003 464
rect 803 400 1003 447
rect 1061 447 1111 464
rect 1211 464 1227 481
rect 1353 481 1485 497
rect 1353 464 1369 481
rect 1211 447 1261 464
rect 1061 400 1261 447
rect 1319 447 1369 464
rect 1469 464 1485 481
rect 1469 447 1519 464
rect 1319 400 1519 447
rect -1519 -447 -1319 -400
rect -1519 -464 -1469 -447
rect -1485 -481 -1469 -464
rect -1369 -464 -1319 -447
rect -1261 -447 -1061 -400
rect -1261 -464 -1211 -447
rect -1369 -481 -1353 -464
rect -1485 -497 -1353 -481
rect -1227 -481 -1211 -464
rect -1111 -464 -1061 -447
rect -1003 -447 -803 -400
rect -1003 -464 -953 -447
rect -1111 -481 -1095 -464
rect -1227 -497 -1095 -481
rect -969 -481 -953 -464
rect -853 -464 -803 -447
rect -745 -447 -545 -400
rect -745 -464 -695 -447
rect -853 -481 -837 -464
rect -969 -497 -837 -481
rect -711 -481 -695 -464
rect -595 -464 -545 -447
rect -487 -447 -287 -400
rect -487 -464 -437 -447
rect -595 -481 -579 -464
rect -711 -497 -579 -481
rect -453 -481 -437 -464
rect -337 -464 -287 -447
rect -229 -447 -29 -400
rect -229 -464 -179 -447
rect -337 -481 -321 -464
rect -453 -497 -321 -481
rect -195 -481 -179 -464
rect -79 -464 -29 -447
rect 29 -447 229 -400
rect 29 -464 79 -447
rect -79 -481 -63 -464
rect -195 -497 -63 -481
rect 63 -481 79 -464
rect 179 -464 229 -447
rect 287 -447 487 -400
rect 287 -464 337 -447
rect 179 -481 195 -464
rect 63 -497 195 -481
rect 321 -481 337 -464
rect 437 -464 487 -447
rect 545 -447 745 -400
rect 545 -464 595 -447
rect 437 -481 453 -464
rect 321 -497 453 -481
rect 579 -481 595 -464
rect 695 -464 745 -447
rect 803 -447 1003 -400
rect 803 -464 853 -447
rect 695 -481 711 -464
rect 579 -497 711 -481
rect 837 -481 853 -464
rect 953 -464 1003 -447
rect 1061 -447 1261 -400
rect 1061 -464 1111 -447
rect 953 -481 969 -464
rect 837 -497 969 -481
rect 1095 -481 1111 -464
rect 1211 -464 1261 -447
rect 1319 -447 1519 -400
rect 1319 -464 1369 -447
rect 1211 -481 1227 -464
rect 1095 -497 1227 -481
rect 1353 -481 1369 -464
rect 1469 -464 1519 -447
rect 1469 -481 1485 -464
rect 1353 -497 1485 -481
<< polycont >>
rect -1469 447 -1369 481
rect -1211 447 -1111 481
rect -953 447 -853 481
rect -695 447 -595 481
rect -437 447 -337 481
rect -179 447 -79 481
rect 79 447 179 481
rect 337 447 437 481
rect 595 447 695 481
rect 853 447 953 481
rect 1111 447 1211 481
rect 1369 447 1469 481
rect -1469 -481 -1369 -447
rect -1211 -481 -1111 -447
rect -953 -481 -853 -447
rect -695 -481 -595 -447
rect -437 -481 -337 -447
rect -179 -481 -79 -447
rect 79 -481 179 -447
rect 337 -481 437 -447
rect 595 -481 695 -447
rect 853 -481 953 -447
rect 1111 -481 1211 -447
rect 1369 -481 1469 -447
<< locali >>
rect -1699 585 -1603 619
rect 1603 585 1699 619
rect -1699 523 -1665 585
rect 1665 523 1699 585
rect -1485 447 -1469 481
rect -1369 447 -1353 481
rect -1227 447 -1211 481
rect -1111 447 -1095 481
rect -969 447 -953 481
rect -853 447 -837 481
rect -711 447 -695 481
rect -595 447 -579 481
rect -453 447 -437 481
rect -337 447 -321 481
rect -195 447 -179 481
rect -79 447 -63 481
rect 63 447 79 481
rect 179 447 195 481
rect 321 447 337 481
rect 437 447 453 481
rect 579 447 595 481
rect 695 447 711 481
rect 837 447 853 481
rect 953 447 969 481
rect 1095 447 1111 481
rect 1211 447 1227 481
rect 1353 447 1369 481
rect 1469 447 1485 481
rect -1565 388 -1531 404
rect -1565 -404 -1531 -388
rect -1307 388 -1273 404
rect -1307 -404 -1273 -388
rect -1049 388 -1015 404
rect -1049 -404 -1015 -388
rect -791 388 -757 404
rect -791 -404 -757 -388
rect -533 388 -499 404
rect -533 -404 -499 -388
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect 499 388 533 404
rect 499 -404 533 -388
rect 757 388 791 404
rect 757 -404 791 -388
rect 1015 388 1049 404
rect 1015 -404 1049 -388
rect 1273 388 1307 404
rect 1273 -404 1307 -388
rect 1531 388 1565 404
rect 1531 -404 1565 -388
rect -1485 -481 -1469 -447
rect -1369 -481 -1353 -447
rect -1227 -481 -1211 -447
rect -1111 -481 -1095 -447
rect -969 -481 -953 -447
rect -853 -481 -837 -447
rect -711 -481 -695 -447
rect -595 -481 -579 -447
rect -453 -481 -437 -447
rect -337 -481 -321 -447
rect -195 -481 -179 -447
rect -79 -481 -63 -447
rect 63 -481 79 -447
rect 179 -481 195 -447
rect 321 -481 337 -447
rect 437 -481 453 -447
rect 579 -481 595 -447
rect 695 -481 711 -447
rect 837 -481 853 -447
rect 953 -481 969 -447
rect 1095 -481 1111 -447
rect 1211 -481 1227 -447
rect 1353 -481 1369 -447
rect 1469 -481 1485 -447
rect -1699 -585 -1665 -523
rect 1665 -585 1699 -523
rect -1699 -619 -1603 -585
rect 1603 -619 1699 -585
<< viali >>
rect -1469 447 -1369 481
rect -1211 447 -1111 481
rect -953 447 -853 481
rect -695 447 -595 481
rect -437 447 -337 481
rect -179 447 -79 481
rect 79 447 179 481
rect 337 447 437 481
rect 595 447 695 481
rect 853 447 953 481
rect 1111 447 1211 481
rect 1369 447 1469 481
rect -1565 -388 -1531 388
rect -1307 -388 -1273 388
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect 1273 -388 1307 388
rect 1531 -388 1565 388
rect -1469 -481 -1369 -447
rect -1211 -481 -1111 -447
rect -953 -481 -853 -447
rect -695 -481 -595 -447
rect -437 -481 -337 -447
rect -179 -481 -79 -447
rect 79 -481 179 -447
rect 337 -481 437 -447
rect 595 -481 695 -447
rect 853 -481 953 -447
rect 1111 -481 1211 -447
rect 1369 -481 1469 -447
<< metal1 >>
rect -1481 481 -1357 487
rect -1481 447 -1469 481
rect -1369 447 -1357 481
rect -1481 441 -1357 447
rect -1223 481 -1099 487
rect -1223 447 -1211 481
rect -1111 447 -1099 481
rect -1223 441 -1099 447
rect -965 481 -841 487
rect -965 447 -953 481
rect -853 447 -841 481
rect -965 441 -841 447
rect -707 481 -583 487
rect -707 447 -695 481
rect -595 447 -583 481
rect -707 441 -583 447
rect -449 481 -325 487
rect -449 447 -437 481
rect -337 447 -325 481
rect -449 441 -325 447
rect -191 481 -67 487
rect -191 447 -179 481
rect -79 447 -67 481
rect -191 441 -67 447
rect 67 481 191 487
rect 67 447 79 481
rect 179 447 191 481
rect 67 441 191 447
rect 325 481 449 487
rect 325 447 337 481
rect 437 447 449 481
rect 325 441 449 447
rect 583 481 707 487
rect 583 447 595 481
rect 695 447 707 481
rect 583 441 707 447
rect 841 481 965 487
rect 841 447 853 481
rect 953 447 965 481
rect 841 441 965 447
rect 1099 481 1223 487
rect 1099 447 1111 481
rect 1211 447 1223 481
rect 1099 441 1223 447
rect 1357 481 1481 487
rect 1357 447 1369 481
rect 1469 447 1481 481
rect 1357 441 1481 447
rect -1571 388 -1525 400
rect -1571 -388 -1565 388
rect -1531 -388 -1525 388
rect -1571 -400 -1525 -388
rect -1313 388 -1267 400
rect -1313 -388 -1307 388
rect -1273 -388 -1267 388
rect -1313 -400 -1267 -388
rect -1055 388 -1009 400
rect -1055 -388 -1049 388
rect -1015 -388 -1009 388
rect -1055 -400 -1009 -388
rect -797 388 -751 400
rect -797 -388 -791 388
rect -757 -388 -751 388
rect -797 -400 -751 -388
rect -539 388 -493 400
rect -539 -388 -533 388
rect -499 -388 -493 388
rect -539 -400 -493 -388
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect 493 388 539 400
rect 493 -388 499 388
rect 533 -388 539 388
rect 493 -400 539 -388
rect 751 388 797 400
rect 751 -388 757 388
rect 791 -388 797 388
rect 751 -400 797 -388
rect 1009 388 1055 400
rect 1009 -388 1015 388
rect 1049 -388 1055 388
rect 1009 -400 1055 -388
rect 1267 388 1313 400
rect 1267 -388 1273 388
rect 1307 -388 1313 388
rect 1267 -400 1313 -388
rect 1525 388 1571 400
rect 1525 -388 1531 388
rect 1565 -388 1571 388
rect 1525 -400 1571 -388
rect -1481 -447 -1357 -441
rect -1481 -481 -1469 -447
rect -1369 -481 -1357 -447
rect -1481 -487 -1357 -481
rect -1223 -447 -1099 -441
rect -1223 -481 -1211 -447
rect -1111 -481 -1099 -447
rect -1223 -487 -1099 -481
rect -965 -447 -841 -441
rect -965 -481 -953 -447
rect -853 -481 -841 -447
rect -965 -487 -841 -481
rect -707 -447 -583 -441
rect -707 -481 -695 -447
rect -595 -481 -583 -447
rect -707 -487 -583 -481
rect -449 -447 -325 -441
rect -449 -481 -437 -447
rect -337 -481 -325 -447
rect -449 -487 -325 -481
rect -191 -447 -67 -441
rect -191 -481 -179 -447
rect -79 -481 -67 -447
rect -191 -487 -67 -481
rect 67 -447 191 -441
rect 67 -481 79 -447
rect 179 -481 191 -447
rect 67 -487 191 -481
rect 325 -447 449 -441
rect 325 -481 337 -447
rect 437 -481 449 -447
rect 325 -487 449 -481
rect 583 -447 707 -441
rect 583 -481 595 -447
rect 695 -481 707 -447
rect 583 -487 707 -481
rect 841 -447 965 -441
rect 841 -481 853 -447
rect 953 -481 965 -447
rect 841 -487 965 -481
rect 1099 -447 1223 -441
rect 1099 -481 1111 -447
rect 1211 -481 1223 -447
rect 1099 -487 1223 -481
rect 1357 -447 1481 -441
rect 1357 -481 1369 -447
rect 1469 -481 1481 -447
rect 1357 -487 1481 -481
<< properties >>
string FIXED_BBOX -1682 -602 1682 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 12 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

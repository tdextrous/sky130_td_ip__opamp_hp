magic
tech sky130A
magscale 1 2
timestamp 1713332875
<< nwell >>
rect -4873 -697 4873 697
<< mvpmos >>
rect -4615 -400 -4415 400
rect -4357 -400 -4157 400
rect -4099 -400 -3899 400
rect -3841 -400 -3641 400
rect -3583 -400 -3383 400
rect -3325 -400 -3125 400
rect -3067 -400 -2867 400
rect -2809 -400 -2609 400
rect -2551 -400 -2351 400
rect -2293 -400 -2093 400
rect -2035 -400 -1835 400
rect -1777 -400 -1577 400
rect -1519 -400 -1319 400
rect -1261 -400 -1061 400
rect -1003 -400 -803 400
rect -745 -400 -545 400
rect -487 -400 -287 400
rect -229 -400 -29 400
rect 29 -400 229 400
rect 287 -400 487 400
rect 545 -400 745 400
rect 803 -400 1003 400
rect 1061 -400 1261 400
rect 1319 -400 1519 400
rect 1577 -400 1777 400
rect 1835 -400 2035 400
rect 2093 -400 2293 400
rect 2351 -400 2551 400
rect 2609 -400 2809 400
rect 2867 -400 3067 400
rect 3125 -400 3325 400
rect 3383 -400 3583 400
rect 3641 -400 3841 400
rect 3899 -400 4099 400
rect 4157 -400 4357 400
rect 4415 -400 4615 400
<< mvpdiff >>
rect -4673 388 -4615 400
rect -4673 -388 -4661 388
rect -4627 -388 -4615 388
rect -4673 -400 -4615 -388
rect -4415 388 -4357 400
rect -4415 -388 -4403 388
rect -4369 -388 -4357 388
rect -4415 -400 -4357 -388
rect -4157 388 -4099 400
rect -4157 -388 -4145 388
rect -4111 -388 -4099 388
rect -4157 -400 -4099 -388
rect -3899 388 -3841 400
rect -3899 -388 -3887 388
rect -3853 -388 -3841 388
rect -3899 -400 -3841 -388
rect -3641 388 -3583 400
rect -3641 -388 -3629 388
rect -3595 -388 -3583 388
rect -3641 -400 -3583 -388
rect -3383 388 -3325 400
rect -3383 -388 -3371 388
rect -3337 -388 -3325 388
rect -3383 -400 -3325 -388
rect -3125 388 -3067 400
rect -3125 -388 -3113 388
rect -3079 -388 -3067 388
rect -3125 -400 -3067 -388
rect -2867 388 -2809 400
rect -2867 -388 -2855 388
rect -2821 -388 -2809 388
rect -2867 -400 -2809 -388
rect -2609 388 -2551 400
rect -2609 -388 -2597 388
rect -2563 -388 -2551 388
rect -2609 -400 -2551 -388
rect -2351 388 -2293 400
rect -2351 -388 -2339 388
rect -2305 -388 -2293 388
rect -2351 -400 -2293 -388
rect -2093 388 -2035 400
rect -2093 -388 -2081 388
rect -2047 -388 -2035 388
rect -2093 -400 -2035 -388
rect -1835 388 -1777 400
rect -1835 -388 -1823 388
rect -1789 -388 -1777 388
rect -1835 -400 -1777 -388
rect -1577 388 -1519 400
rect -1577 -388 -1565 388
rect -1531 -388 -1519 388
rect -1577 -400 -1519 -388
rect -1319 388 -1261 400
rect -1319 -388 -1307 388
rect -1273 -388 -1261 388
rect -1319 -400 -1261 -388
rect -1061 388 -1003 400
rect -1061 -388 -1049 388
rect -1015 -388 -1003 388
rect -1061 -400 -1003 -388
rect -803 388 -745 400
rect -803 -388 -791 388
rect -757 -388 -745 388
rect -803 -400 -745 -388
rect -545 388 -487 400
rect -545 -388 -533 388
rect -499 -388 -487 388
rect -545 -400 -487 -388
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect 487 388 545 400
rect 487 -388 499 388
rect 533 -388 545 388
rect 487 -400 545 -388
rect 745 388 803 400
rect 745 -388 757 388
rect 791 -388 803 388
rect 745 -400 803 -388
rect 1003 388 1061 400
rect 1003 -388 1015 388
rect 1049 -388 1061 388
rect 1003 -400 1061 -388
rect 1261 388 1319 400
rect 1261 -388 1273 388
rect 1307 -388 1319 388
rect 1261 -400 1319 -388
rect 1519 388 1577 400
rect 1519 -388 1531 388
rect 1565 -388 1577 388
rect 1519 -400 1577 -388
rect 1777 388 1835 400
rect 1777 -388 1789 388
rect 1823 -388 1835 388
rect 1777 -400 1835 -388
rect 2035 388 2093 400
rect 2035 -388 2047 388
rect 2081 -388 2093 388
rect 2035 -400 2093 -388
rect 2293 388 2351 400
rect 2293 -388 2305 388
rect 2339 -388 2351 388
rect 2293 -400 2351 -388
rect 2551 388 2609 400
rect 2551 -388 2563 388
rect 2597 -388 2609 388
rect 2551 -400 2609 -388
rect 2809 388 2867 400
rect 2809 -388 2821 388
rect 2855 -388 2867 388
rect 2809 -400 2867 -388
rect 3067 388 3125 400
rect 3067 -388 3079 388
rect 3113 -388 3125 388
rect 3067 -400 3125 -388
rect 3325 388 3383 400
rect 3325 -388 3337 388
rect 3371 -388 3383 388
rect 3325 -400 3383 -388
rect 3583 388 3641 400
rect 3583 -388 3595 388
rect 3629 -388 3641 388
rect 3583 -400 3641 -388
rect 3841 388 3899 400
rect 3841 -388 3853 388
rect 3887 -388 3899 388
rect 3841 -400 3899 -388
rect 4099 388 4157 400
rect 4099 -388 4111 388
rect 4145 -388 4157 388
rect 4099 -400 4157 -388
rect 4357 388 4415 400
rect 4357 -388 4369 388
rect 4403 -388 4415 388
rect 4357 -400 4415 -388
rect 4615 388 4673 400
rect 4615 -388 4627 388
rect 4661 -388 4673 388
rect 4615 -400 4673 -388
<< mvpdiffc >>
rect -4661 -388 -4627 388
rect -4403 -388 -4369 388
rect -4145 -388 -4111 388
rect -3887 -388 -3853 388
rect -3629 -388 -3595 388
rect -3371 -388 -3337 388
rect -3113 -388 -3079 388
rect -2855 -388 -2821 388
rect -2597 -388 -2563 388
rect -2339 -388 -2305 388
rect -2081 -388 -2047 388
rect -1823 -388 -1789 388
rect -1565 -388 -1531 388
rect -1307 -388 -1273 388
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect 1273 -388 1307 388
rect 1531 -388 1565 388
rect 1789 -388 1823 388
rect 2047 -388 2081 388
rect 2305 -388 2339 388
rect 2563 -388 2597 388
rect 2821 -388 2855 388
rect 3079 -388 3113 388
rect 3337 -388 3371 388
rect 3595 -388 3629 388
rect 3853 -388 3887 388
rect 4111 -388 4145 388
rect 4369 -388 4403 388
rect 4627 -388 4661 388
<< mvnsubdiff >>
rect -4807 619 4807 631
rect -4807 585 -4699 619
rect 4699 585 4807 619
rect -4807 573 4807 585
rect -4807 523 -4749 573
rect -4807 -523 -4795 523
rect -4761 -523 -4749 523
rect 4749 523 4807 573
rect -4807 -573 -4749 -523
rect 4749 -523 4761 523
rect 4795 -523 4807 523
rect 4749 -573 4807 -523
rect -4807 -585 4807 -573
rect -4807 -619 -4699 -585
rect 4699 -619 4807 -585
rect -4807 -631 4807 -619
<< mvnsubdiffcont >>
rect -4699 585 4699 619
rect -4795 -523 -4761 523
rect 4761 -523 4795 523
rect -4699 -619 4699 -585
<< poly >>
rect -4581 481 -4449 497
rect -4581 464 -4565 481
rect -4615 447 -4565 464
rect -4465 464 -4449 481
rect -4323 481 -4191 497
rect -4323 464 -4307 481
rect -4465 447 -4415 464
rect -4615 400 -4415 447
rect -4357 447 -4307 464
rect -4207 464 -4191 481
rect -4065 481 -3933 497
rect -4065 464 -4049 481
rect -4207 447 -4157 464
rect -4357 400 -4157 447
rect -4099 447 -4049 464
rect -3949 464 -3933 481
rect -3807 481 -3675 497
rect -3807 464 -3791 481
rect -3949 447 -3899 464
rect -4099 400 -3899 447
rect -3841 447 -3791 464
rect -3691 464 -3675 481
rect -3549 481 -3417 497
rect -3549 464 -3533 481
rect -3691 447 -3641 464
rect -3841 400 -3641 447
rect -3583 447 -3533 464
rect -3433 464 -3417 481
rect -3291 481 -3159 497
rect -3291 464 -3275 481
rect -3433 447 -3383 464
rect -3583 400 -3383 447
rect -3325 447 -3275 464
rect -3175 464 -3159 481
rect -3033 481 -2901 497
rect -3033 464 -3017 481
rect -3175 447 -3125 464
rect -3325 400 -3125 447
rect -3067 447 -3017 464
rect -2917 464 -2901 481
rect -2775 481 -2643 497
rect -2775 464 -2759 481
rect -2917 447 -2867 464
rect -3067 400 -2867 447
rect -2809 447 -2759 464
rect -2659 464 -2643 481
rect -2517 481 -2385 497
rect -2517 464 -2501 481
rect -2659 447 -2609 464
rect -2809 400 -2609 447
rect -2551 447 -2501 464
rect -2401 464 -2385 481
rect -2259 481 -2127 497
rect -2259 464 -2243 481
rect -2401 447 -2351 464
rect -2551 400 -2351 447
rect -2293 447 -2243 464
rect -2143 464 -2127 481
rect -2001 481 -1869 497
rect -2001 464 -1985 481
rect -2143 447 -2093 464
rect -2293 400 -2093 447
rect -2035 447 -1985 464
rect -1885 464 -1869 481
rect -1743 481 -1611 497
rect -1743 464 -1727 481
rect -1885 447 -1835 464
rect -2035 400 -1835 447
rect -1777 447 -1727 464
rect -1627 464 -1611 481
rect -1485 481 -1353 497
rect -1485 464 -1469 481
rect -1627 447 -1577 464
rect -1777 400 -1577 447
rect -1519 447 -1469 464
rect -1369 464 -1353 481
rect -1227 481 -1095 497
rect -1227 464 -1211 481
rect -1369 447 -1319 464
rect -1519 400 -1319 447
rect -1261 447 -1211 464
rect -1111 464 -1095 481
rect -969 481 -837 497
rect -969 464 -953 481
rect -1111 447 -1061 464
rect -1261 400 -1061 447
rect -1003 447 -953 464
rect -853 464 -837 481
rect -711 481 -579 497
rect -711 464 -695 481
rect -853 447 -803 464
rect -1003 400 -803 447
rect -745 447 -695 464
rect -595 464 -579 481
rect -453 481 -321 497
rect -453 464 -437 481
rect -595 447 -545 464
rect -745 400 -545 447
rect -487 447 -437 464
rect -337 464 -321 481
rect -195 481 -63 497
rect -195 464 -179 481
rect -337 447 -287 464
rect -487 400 -287 447
rect -229 447 -179 464
rect -79 464 -63 481
rect 63 481 195 497
rect 63 464 79 481
rect -79 447 -29 464
rect -229 400 -29 447
rect 29 447 79 464
rect 179 464 195 481
rect 321 481 453 497
rect 321 464 337 481
rect 179 447 229 464
rect 29 400 229 447
rect 287 447 337 464
rect 437 464 453 481
rect 579 481 711 497
rect 579 464 595 481
rect 437 447 487 464
rect 287 400 487 447
rect 545 447 595 464
rect 695 464 711 481
rect 837 481 969 497
rect 837 464 853 481
rect 695 447 745 464
rect 545 400 745 447
rect 803 447 853 464
rect 953 464 969 481
rect 1095 481 1227 497
rect 1095 464 1111 481
rect 953 447 1003 464
rect 803 400 1003 447
rect 1061 447 1111 464
rect 1211 464 1227 481
rect 1353 481 1485 497
rect 1353 464 1369 481
rect 1211 447 1261 464
rect 1061 400 1261 447
rect 1319 447 1369 464
rect 1469 464 1485 481
rect 1611 481 1743 497
rect 1611 464 1627 481
rect 1469 447 1519 464
rect 1319 400 1519 447
rect 1577 447 1627 464
rect 1727 464 1743 481
rect 1869 481 2001 497
rect 1869 464 1885 481
rect 1727 447 1777 464
rect 1577 400 1777 447
rect 1835 447 1885 464
rect 1985 464 2001 481
rect 2127 481 2259 497
rect 2127 464 2143 481
rect 1985 447 2035 464
rect 1835 400 2035 447
rect 2093 447 2143 464
rect 2243 464 2259 481
rect 2385 481 2517 497
rect 2385 464 2401 481
rect 2243 447 2293 464
rect 2093 400 2293 447
rect 2351 447 2401 464
rect 2501 464 2517 481
rect 2643 481 2775 497
rect 2643 464 2659 481
rect 2501 447 2551 464
rect 2351 400 2551 447
rect 2609 447 2659 464
rect 2759 464 2775 481
rect 2901 481 3033 497
rect 2901 464 2917 481
rect 2759 447 2809 464
rect 2609 400 2809 447
rect 2867 447 2917 464
rect 3017 464 3033 481
rect 3159 481 3291 497
rect 3159 464 3175 481
rect 3017 447 3067 464
rect 2867 400 3067 447
rect 3125 447 3175 464
rect 3275 464 3291 481
rect 3417 481 3549 497
rect 3417 464 3433 481
rect 3275 447 3325 464
rect 3125 400 3325 447
rect 3383 447 3433 464
rect 3533 464 3549 481
rect 3675 481 3807 497
rect 3675 464 3691 481
rect 3533 447 3583 464
rect 3383 400 3583 447
rect 3641 447 3691 464
rect 3791 464 3807 481
rect 3933 481 4065 497
rect 3933 464 3949 481
rect 3791 447 3841 464
rect 3641 400 3841 447
rect 3899 447 3949 464
rect 4049 464 4065 481
rect 4191 481 4323 497
rect 4191 464 4207 481
rect 4049 447 4099 464
rect 3899 400 4099 447
rect 4157 447 4207 464
rect 4307 464 4323 481
rect 4449 481 4581 497
rect 4449 464 4465 481
rect 4307 447 4357 464
rect 4157 400 4357 447
rect 4415 447 4465 464
rect 4565 464 4581 481
rect 4565 447 4615 464
rect 4415 400 4615 447
rect -4615 -447 -4415 -400
rect -4615 -464 -4565 -447
rect -4581 -481 -4565 -464
rect -4465 -464 -4415 -447
rect -4357 -447 -4157 -400
rect -4357 -464 -4307 -447
rect -4465 -481 -4449 -464
rect -4581 -497 -4449 -481
rect -4323 -481 -4307 -464
rect -4207 -464 -4157 -447
rect -4099 -447 -3899 -400
rect -4099 -464 -4049 -447
rect -4207 -481 -4191 -464
rect -4323 -497 -4191 -481
rect -4065 -481 -4049 -464
rect -3949 -464 -3899 -447
rect -3841 -447 -3641 -400
rect -3841 -464 -3791 -447
rect -3949 -481 -3933 -464
rect -4065 -497 -3933 -481
rect -3807 -481 -3791 -464
rect -3691 -464 -3641 -447
rect -3583 -447 -3383 -400
rect -3583 -464 -3533 -447
rect -3691 -481 -3675 -464
rect -3807 -497 -3675 -481
rect -3549 -481 -3533 -464
rect -3433 -464 -3383 -447
rect -3325 -447 -3125 -400
rect -3325 -464 -3275 -447
rect -3433 -481 -3417 -464
rect -3549 -497 -3417 -481
rect -3291 -481 -3275 -464
rect -3175 -464 -3125 -447
rect -3067 -447 -2867 -400
rect -3067 -464 -3017 -447
rect -3175 -481 -3159 -464
rect -3291 -497 -3159 -481
rect -3033 -481 -3017 -464
rect -2917 -464 -2867 -447
rect -2809 -447 -2609 -400
rect -2809 -464 -2759 -447
rect -2917 -481 -2901 -464
rect -3033 -497 -2901 -481
rect -2775 -481 -2759 -464
rect -2659 -464 -2609 -447
rect -2551 -447 -2351 -400
rect -2551 -464 -2501 -447
rect -2659 -481 -2643 -464
rect -2775 -497 -2643 -481
rect -2517 -481 -2501 -464
rect -2401 -464 -2351 -447
rect -2293 -447 -2093 -400
rect -2293 -464 -2243 -447
rect -2401 -481 -2385 -464
rect -2517 -497 -2385 -481
rect -2259 -481 -2243 -464
rect -2143 -464 -2093 -447
rect -2035 -447 -1835 -400
rect -2035 -464 -1985 -447
rect -2143 -481 -2127 -464
rect -2259 -497 -2127 -481
rect -2001 -481 -1985 -464
rect -1885 -464 -1835 -447
rect -1777 -447 -1577 -400
rect -1777 -464 -1727 -447
rect -1885 -481 -1869 -464
rect -2001 -497 -1869 -481
rect -1743 -481 -1727 -464
rect -1627 -464 -1577 -447
rect -1519 -447 -1319 -400
rect -1519 -464 -1469 -447
rect -1627 -481 -1611 -464
rect -1743 -497 -1611 -481
rect -1485 -481 -1469 -464
rect -1369 -464 -1319 -447
rect -1261 -447 -1061 -400
rect -1261 -464 -1211 -447
rect -1369 -481 -1353 -464
rect -1485 -497 -1353 -481
rect -1227 -481 -1211 -464
rect -1111 -464 -1061 -447
rect -1003 -447 -803 -400
rect -1003 -464 -953 -447
rect -1111 -481 -1095 -464
rect -1227 -497 -1095 -481
rect -969 -481 -953 -464
rect -853 -464 -803 -447
rect -745 -447 -545 -400
rect -745 -464 -695 -447
rect -853 -481 -837 -464
rect -969 -497 -837 -481
rect -711 -481 -695 -464
rect -595 -464 -545 -447
rect -487 -447 -287 -400
rect -487 -464 -437 -447
rect -595 -481 -579 -464
rect -711 -497 -579 -481
rect -453 -481 -437 -464
rect -337 -464 -287 -447
rect -229 -447 -29 -400
rect -229 -464 -179 -447
rect -337 -481 -321 -464
rect -453 -497 -321 -481
rect -195 -481 -179 -464
rect -79 -464 -29 -447
rect 29 -447 229 -400
rect 29 -464 79 -447
rect -79 -481 -63 -464
rect -195 -497 -63 -481
rect 63 -481 79 -464
rect 179 -464 229 -447
rect 287 -447 487 -400
rect 287 -464 337 -447
rect 179 -481 195 -464
rect 63 -497 195 -481
rect 321 -481 337 -464
rect 437 -464 487 -447
rect 545 -447 745 -400
rect 545 -464 595 -447
rect 437 -481 453 -464
rect 321 -497 453 -481
rect 579 -481 595 -464
rect 695 -464 745 -447
rect 803 -447 1003 -400
rect 803 -464 853 -447
rect 695 -481 711 -464
rect 579 -497 711 -481
rect 837 -481 853 -464
rect 953 -464 1003 -447
rect 1061 -447 1261 -400
rect 1061 -464 1111 -447
rect 953 -481 969 -464
rect 837 -497 969 -481
rect 1095 -481 1111 -464
rect 1211 -464 1261 -447
rect 1319 -447 1519 -400
rect 1319 -464 1369 -447
rect 1211 -481 1227 -464
rect 1095 -497 1227 -481
rect 1353 -481 1369 -464
rect 1469 -464 1519 -447
rect 1577 -447 1777 -400
rect 1577 -464 1627 -447
rect 1469 -481 1485 -464
rect 1353 -497 1485 -481
rect 1611 -481 1627 -464
rect 1727 -464 1777 -447
rect 1835 -447 2035 -400
rect 1835 -464 1885 -447
rect 1727 -481 1743 -464
rect 1611 -497 1743 -481
rect 1869 -481 1885 -464
rect 1985 -464 2035 -447
rect 2093 -447 2293 -400
rect 2093 -464 2143 -447
rect 1985 -481 2001 -464
rect 1869 -497 2001 -481
rect 2127 -481 2143 -464
rect 2243 -464 2293 -447
rect 2351 -447 2551 -400
rect 2351 -464 2401 -447
rect 2243 -481 2259 -464
rect 2127 -497 2259 -481
rect 2385 -481 2401 -464
rect 2501 -464 2551 -447
rect 2609 -447 2809 -400
rect 2609 -464 2659 -447
rect 2501 -481 2517 -464
rect 2385 -497 2517 -481
rect 2643 -481 2659 -464
rect 2759 -464 2809 -447
rect 2867 -447 3067 -400
rect 2867 -464 2917 -447
rect 2759 -481 2775 -464
rect 2643 -497 2775 -481
rect 2901 -481 2917 -464
rect 3017 -464 3067 -447
rect 3125 -447 3325 -400
rect 3125 -464 3175 -447
rect 3017 -481 3033 -464
rect 2901 -497 3033 -481
rect 3159 -481 3175 -464
rect 3275 -464 3325 -447
rect 3383 -447 3583 -400
rect 3383 -464 3433 -447
rect 3275 -481 3291 -464
rect 3159 -497 3291 -481
rect 3417 -481 3433 -464
rect 3533 -464 3583 -447
rect 3641 -447 3841 -400
rect 3641 -464 3691 -447
rect 3533 -481 3549 -464
rect 3417 -497 3549 -481
rect 3675 -481 3691 -464
rect 3791 -464 3841 -447
rect 3899 -447 4099 -400
rect 3899 -464 3949 -447
rect 3791 -481 3807 -464
rect 3675 -497 3807 -481
rect 3933 -481 3949 -464
rect 4049 -464 4099 -447
rect 4157 -447 4357 -400
rect 4157 -464 4207 -447
rect 4049 -481 4065 -464
rect 3933 -497 4065 -481
rect 4191 -481 4207 -464
rect 4307 -464 4357 -447
rect 4415 -447 4615 -400
rect 4415 -464 4465 -447
rect 4307 -481 4323 -464
rect 4191 -497 4323 -481
rect 4449 -481 4465 -464
rect 4565 -464 4615 -447
rect 4565 -481 4581 -464
rect 4449 -497 4581 -481
<< polycont >>
rect -4565 447 -4465 481
rect -4307 447 -4207 481
rect -4049 447 -3949 481
rect -3791 447 -3691 481
rect -3533 447 -3433 481
rect -3275 447 -3175 481
rect -3017 447 -2917 481
rect -2759 447 -2659 481
rect -2501 447 -2401 481
rect -2243 447 -2143 481
rect -1985 447 -1885 481
rect -1727 447 -1627 481
rect -1469 447 -1369 481
rect -1211 447 -1111 481
rect -953 447 -853 481
rect -695 447 -595 481
rect -437 447 -337 481
rect -179 447 -79 481
rect 79 447 179 481
rect 337 447 437 481
rect 595 447 695 481
rect 853 447 953 481
rect 1111 447 1211 481
rect 1369 447 1469 481
rect 1627 447 1727 481
rect 1885 447 1985 481
rect 2143 447 2243 481
rect 2401 447 2501 481
rect 2659 447 2759 481
rect 2917 447 3017 481
rect 3175 447 3275 481
rect 3433 447 3533 481
rect 3691 447 3791 481
rect 3949 447 4049 481
rect 4207 447 4307 481
rect 4465 447 4565 481
rect -4565 -481 -4465 -447
rect -4307 -481 -4207 -447
rect -4049 -481 -3949 -447
rect -3791 -481 -3691 -447
rect -3533 -481 -3433 -447
rect -3275 -481 -3175 -447
rect -3017 -481 -2917 -447
rect -2759 -481 -2659 -447
rect -2501 -481 -2401 -447
rect -2243 -481 -2143 -447
rect -1985 -481 -1885 -447
rect -1727 -481 -1627 -447
rect -1469 -481 -1369 -447
rect -1211 -481 -1111 -447
rect -953 -481 -853 -447
rect -695 -481 -595 -447
rect -437 -481 -337 -447
rect -179 -481 -79 -447
rect 79 -481 179 -447
rect 337 -481 437 -447
rect 595 -481 695 -447
rect 853 -481 953 -447
rect 1111 -481 1211 -447
rect 1369 -481 1469 -447
rect 1627 -481 1727 -447
rect 1885 -481 1985 -447
rect 2143 -481 2243 -447
rect 2401 -481 2501 -447
rect 2659 -481 2759 -447
rect 2917 -481 3017 -447
rect 3175 -481 3275 -447
rect 3433 -481 3533 -447
rect 3691 -481 3791 -447
rect 3949 -481 4049 -447
rect 4207 -481 4307 -447
rect 4465 -481 4565 -447
<< locali >>
rect -4795 585 -4699 619
rect 4699 585 4795 619
rect -4795 523 -4761 585
rect 4761 523 4795 585
rect -4581 447 -4565 481
rect -4465 447 -4449 481
rect -4323 447 -4307 481
rect -4207 447 -4191 481
rect -4065 447 -4049 481
rect -3949 447 -3933 481
rect -3807 447 -3791 481
rect -3691 447 -3675 481
rect -3549 447 -3533 481
rect -3433 447 -3417 481
rect -3291 447 -3275 481
rect -3175 447 -3159 481
rect -3033 447 -3017 481
rect -2917 447 -2901 481
rect -2775 447 -2759 481
rect -2659 447 -2643 481
rect -2517 447 -2501 481
rect -2401 447 -2385 481
rect -2259 447 -2243 481
rect -2143 447 -2127 481
rect -2001 447 -1985 481
rect -1885 447 -1869 481
rect -1743 447 -1727 481
rect -1627 447 -1611 481
rect -1485 447 -1469 481
rect -1369 447 -1353 481
rect -1227 447 -1211 481
rect -1111 447 -1095 481
rect -969 447 -953 481
rect -853 447 -837 481
rect -711 447 -695 481
rect -595 447 -579 481
rect -453 447 -437 481
rect -337 447 -321 481
rect -195 447 -179 481
rect -79 447 -63 481
rect 63 447 79 481
rect 179 447 195 481
rect 321 447 337 481
rect 437 447 453 481
rect 579 447 595 481
rect 695 447 711 481
rect 837 447 853 481
rect 953 447 969 481
rect 1095 447 1111 481
rect 1211 447 1227 481
rect 1353 447 1369 481
rect 1469 447 1485 481
rect 1611 447 1627 481
rect 1727 447 1743 481
rect 1869 447 1885 481
rect 1985 447 2001 481
rect 2127 447 2143 481
rect 2243 447 2259 481
rect 2385 447 2401 481
rect 2501 447 2517 481
rect 2643 447 2659 481
rect 2759 447 2775 481
rect 2901 447 2917 481
rect 3017 447 3033 481
rect 3159 447 3175 481
rect 3275 447 3291 481
rect 3417 447 3433 481
rect 3533 447 3549 481
rect 3675 447 3691 481
rect 3791 447 3807 481
rect 3933 447 3949 481
rect 4049 447 4065 481
rect 4191 447 4207 481
rect 4307 447 4323 481
rect 4449 447 4465 481
rect 4565 447 4581 481
rect -4661 388 -4627 404
rect -4661 -404 -4627 -388
rect -4403 388 -4369 404
rect -4403 -404 -4369 -388
rect -4145 388 -4111 404
rect -4145 -404 -4111 -388
rect -3887 388 -3853 404
rect -3887 -404 -3853 -388
rect -3629 388 -3595 404
rect -3629 -404 -3595 -388
rect -3371 388 -3337 404
rect -3371 -404 -3337 -388
rect -3113 388 -3079 404
rect -3113 -404 -3079 -388
rect -2855 388 -2821 404
rect -2855 -404 -2821 -388
rect -2597 388 -2563 404
rect -2597 -404 -2563 -388
rect -2339 388 -2305 404
rect -2339 -404 -2305 -388
rect -2081 388 -2047 404
rect -2081 -404 -2047 -388
rect -1823 388 -1789 404
rect -1823 -404 -1789 -388
rect -1565 388 -1531 404
rect -1565 -404 -1531 -388
rect -1307 388 -1273 404
rect -1307 -404 -1273 -388
rect -1049 388 -1015 404
rect -1049 -404 -1015 -388
rect -791 388 -757 404
rect -791 -404 -757 -388
rect -533 388 -499 404
rect -533 -404 -499 -388
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect 499 388 533 404
rect 499 -404 533 -388
rect 757 388 791 404
rect 757 -404 791 -388
rect 1015 388 1049 404
rect 1015 -404 1049 -388
rect 1273 388 1307 404
rect 1273 -404 1307 -388
rect 1531 388 1565 404
rect 1531 -404 1565 -388
rect 1789 388 1823 404
rect 1789 -404 1823 -388
rect 2047 388 2081 404
rect 2047 -404 2081 -388
rect 2305 388 2339 404
rect 2305 -404 2339 -388
rect 2563 388 2597 404
rect 2563 -404 2597 -388
rect 2821 388 2855 404
rect 2821 -404 2855 -388
rect 3079 388 3113 404
rect 3079 -404 3113 -388
rect 3337 388 3371 404
rect 3337 -404 3371 -388
rect 3595 388 3629 404
rect 3595 -404 3629 -388
rect 3853 388 3887 404
rect 3853 -404 3887 -388
rect 4111 388 4145 404
rect 4111 -404 4145 -388
rect 4369 388 4403 404
rect 4369 -404 4403 -388
rect 4627 388 4661 404
rect 4627 -404 4661 -388
rect -4581 -481 -4565 -447
rect -4465 -481 -4449 -447
rect -4323 -481 -4307 -447
rect -4207 -481 -4191 -447
rect -4065 -481 -4049 -447
rect -3949 -481 -3933 -447
rect -3807 -481 -3791 -447
rect -3691 -481 -3675 -447
rect -3549 -481 -3533 -447
rect -3433 -481 -3417 -447
rect -3291 -481 -3275 -447
rect -3175 -481 -3159 -447
rect -3033 -481 -3017 -447
rect -2917 -481 -2901 -447
rect -2775 -481 -2759 -447
rect -2659 -481 -2643 -447
rect -2517 -481 -2501 -447
rect -2401 -481 -2385 -447
rect -2259 -481 -2243 -447
rect -2143 -481 -2127 -447
rect -2001 -481 -1985 -447
rect -1885 -481 -1869 -447
rect -1743 -481 -1727 -447
rect -1627 -481 -1611 -447
rect -1485 -481 -1469 -447
rect -1369 -481 -1353 -447
rect -1227 -481 -1211 -447
rect -1111 -481 -1095 -447
rect -969 -481 -953 -447
rect -853 -481 -837 -447
rect -711 -481 -695 -447
rect -595 -481 -579 -447
rect -453 -481 -437 -447
rect -337 -481 -321 -447
rect -195 -481 -179 -447
rect -79 -481 -63 -447
rect 63 -481 79 -447
rect 179 -481 195 -447
rect 321 -481 337 -447
rect 437 -481 453 -447
rect 579 -481 595 -447
rect 695 -481 711 -447
rect 837 -481 853 -447
rect 953 -481 969 -447
rect 1095 -481 1111 -447
rect 1211 -481 1227 -447
rect 1353 -481 1369 -447
rect 1469 -481 1485 -447
rect 1611 -481 1627 -447
rect 1727 -481 1743 -447
rect 1869 -481 1885 -447
rect 1985 -481 2001 -447
rect 2127 -481 2143 -447
rect 2243 -481 2259 -447
rect 2385 -481 2401 -447
rect 2501 -481 2517 -447
rect 2643 -481 2659 -447
rect 2759 -481 2775 -447
rect 2901 -481 2917 -447
rect 3017 -481 3033 -447
rect 3159 -481 3175 -447
rect 3275 -481 3291 -447
rect 3417 -481 3433 -447
rect 3533 -481 3549 -447
rect 3675 -481 3691 -447
rect 3791 -481 3807 -447
rect 3933 -481 3949 -447
rect 4049 -481 4065 -447
rect 4191 -481 4207 -447
rect 4307 -481 4323 -447
rect 4449 -481 4465 -447
rect 4565 -481 4581 -447
rect -4795 -585 -4761 -523
rect 4761 -585 4795 -523
rect -4795 -619 -4699 -585
rect 4699 -619 4795 -585
<< viali >>
rect -4565 447 -4465 481
rect -4307 447 -4207 481
rect -4049 447 -3949 481
rect -3791 447 -3691 481
rect -3533 447 -3433 481
rect -3275 447 -3175 481
rect -3017 447 -2917 481
rect -2759 447 -2659 481
rect -2501 447 -2401 481
rect -2243 447 -2143 481
rect -1985 447 -1885 481
rect -1727 447 -1627 481
rect -1469 447 -1369 481
rect -1211 447 -1111 481
rect -953 447 -853 481
rect -695 447 -595 481
rect -437 447 -337 481
rect -179 447 -79 481
rect 79 447 179 481
rect 337 447 437 481
rect 595 447 695 481
rect 853 447 953 481
rect 1111 447 1211 481
rect 1369 447 1469 481
rect 1627 447 1727 481
rect 1885 447 1985 481
rect 2143 447 2243 481
rect 2401 447 2501 481
rect 2659 447 2759 481
rect 2917 447 3017 481
rect 3175 447 3275 481
rect 3433 447 3533 481
rect 3691 447 3791 481
rect 3949 447 4049 481
rect 4207 447 4307 481
rect 4465 447 4565 481
rect -4661 -388 -4627 388
rect -4403 -388 -4369 388
rect -4145 -388 -4111 388
rect -3887 -388 -3853 388
rect -3629 -388 -3595 388
rect -3371 -388 -3337 388
rect -3113 -388 -3079 388
rect -2855 -388 -2821 388
rect -2597 -388 -2563 388
rect -2339 -388 -2305 388
rect -2081 -388 -2047 388
rect -1823 -388 -1789 388
rect -1565 -388 -1531 388
rect -1307 -388 -1273 388
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect 1273 -388 1307 388
rect 1531 -388 1565 388
rect 1789 -388 1823 388
rect 2047 -388 2081 388
rect 2305 -388 2339 388
rect 2563 -388 2597 388
rect 2821 -388 2855 388
rect 3079 -388 3113 388
rect 3337 -388 3371 388
rect 3595 -388 3629 388
rect 3853 -388 3887 388
rect 4111 -388 4145 388
rect 4369 -388 4403 388
rect 4627 -388 4661 388
rect -4565 -481 -4465 -447
rect -4307 -481 -4207 -447
rect -4049 -481 -3949 -447
rect -3791 -481 -3691 -447
rect -3533 -481 -3433 -447
rect -3275 -481 -3175 -447
rect -3017 -481 -2917 -447
rect -2759 -481 -2659 -447
rect -2501 -481 -2401 -447
rect -2243 -481 -2143 -447
rect -1985 -481 -1885 -447
rect -1727 -481 -1627 -447
rect -1469 -481 -1369 -447
rect -1211 -481 -1111 -447
rect -953 -481 -853 -447
rect -695 -481 -595 -447
rect -437 -481 -337 -447
rect -179 -481 -79 -447
rect 79 -481 179 -447
rect 337 -481 437 -447
rect 595 -481 695 -447
rect 853 -481 953 -447
rect 1111 -481 1211 -447
rect 1369 -481 1469 -447
rect 1627 -481 1727 -447
rect 1885 -481 1985 -447
rect 2143 -481 2243 -447
rect 2401 -481 2501 -447
rect 2659 -481 2759 -447
rect 2917 -481 3017 -447
rect 3175 -481 3275 -447
rect 3433 -481 3533 -447
rect 3691 -481 3791 -447
rect 3949 -481 4049 -447
rect 4207 -481 4307 -447
rect 4465 -481 4565 -447
<< metal1 >>
rect -4577 481 -4453 487
rect -4577 447 -4565 481
rect -4465 447 -4453 481
rect -4577 441 -4453 447
rect -4319 481 -4195 487
rect -4319 447 -4307 481
rect -4207 447 -4195 481
rect -4319 441 -4195 447
rect -4061 481 -3937 487
rect -4061 447 -4049 481
rect -3949 447 -3937 481
rect -4061 441 -3937 447
rect -3803 481 -3679 487
rect -3803 447 -3791 481
rect -3691 447 -3679 481
rect -3803 441 -3679 447
rect -3545 481 -3421 487
rect -3545 447 -3533 481
rect -3433 447 -3421 481
rect -3545 441 -3421 447
rect -3287 481 -3163 487
rect -3287 447 -3275 481
rect -3175 447 -3163 481
rect -3287 441 -3163 447
rect -3029 481 -2905 487
rect -3029 447 -3017 481
rect -2917 447 -2905 481
rect -3029 441 -2905 447
rect -2771 481 -2647 487
rect -2771 447 -2759 481
rect -2659 447 -2647 481
rect -2771 441 -2647 447
rect -2513 481 -2389 487
rect -2513 447 -2501 481
rect -2401 447 -2389 481
rect -2513 441 -2389 447
rect -2255 481 -2131 487
rect -2255 447 -2243 481
rect -2143 447 -2131 481
rect -2255 441 -2131 447
rect -1997 481 -1873 487
rect -1997 447 -1985 481
rect -1885 447 -1873 481
rect -1997 441 -1873 447
rect -1739 481 -1615 487
rect -1739 447 -1727 481
rect -1627 447 -1615 481
rect -1739 441 -1615 447
rect -1481 481 -1357 487
rect -1481 447 -1469 481
rect -1369 447 -1357 481
rect -1481 441 -1357 447
rect -1223 481 -1099 487
rect -1223 447 -1211 481
rect -1111 447 -1099 481
rect -1223 441 -1099 447
rect -965 481 -841 487
rect -965 447 -953 481
rect -853 447 -841 481
rect -965 441 -841 447
rect -707 481 -583 487
rect -707 447 -695 481
rect -595 447 -583 481
rect -707 441 -583 447
rect -449 481 -325 487
rect -449 447 -437 481
rect -337 447 -325 481
rect -449 441 -325 447
rect -191 481 -67 487
rect -191 447 -179 481
rect -79 447 -67 481
rect -191 441 -67 447
rect 67 481 191 487
rect 67 447 79 481
rect 179 447 191 481
rect 67 441 191 447
rect 325 481 449 487
rect 325 447 337 481
rect 437 447 449 481
rect 325 441 449 447
rect 583 481 707 487
rect 583 447 595 481
rect 695 447 707 481
rect 583 441 707 447
rect 841 481 965 487
rect 841 447 853 481
rect 953 447 965 481
rect 841 441 965 447
rect 1099 481 1223 487
rect 1099 447 1111 481
rect 1211 447 1223 481
rect 1099 441 1223 447
rect 1357 481 1481 487
rect 1357 447 1369 481
rect 1469 447 1481 481
rect 1357 441 1481 447
rect 1615 481 1739 487
rect 1615 447 1627 481
rect 1727 447 1739 481
rect 1615 441 1739 447
rect 1873 481 1997 487
rect 1873 447 1885 481
rect 1985 447 1997 481
rect 1873 441 1997 447
rect 2131 481 2255 487
rect 2131 447 2143 481
rect 2243 447 2255 481
rect 2131 441 2255 447
rect 2389 481 2513 487
rect 2389 447 2401 481
rect 2501 447 2513 481
rect 2389 441 2513 447
rect 2647 481 2771 487
rect 2647 447 2659 481
rect 2759 447 2771 481
rect 2647 441 2771 447
rect 2905 481 3029 487
rect 2905 447 2917 481
rect 3017 447 3029 481
rect 2905 441 3029 447
rect 3163 481 3287 487
rect 3163 447 3175 481
rect 3275 447 3287 481
rect 3163 441 3287 447
rect 3421 481 3545 487
rect 3421 447 3433 481
rect 3533 447 3545 481
rect 3421 441 3545 447
rect 3679 481 3803 487
rect 3679 447 3691 481
rect 3791 447 3803 481
rect 3679 441 3803 447
rect 3937 481 4061 487
rect 3937 447 3949 481
rect 4049 447 4061 481
rect 3937 441 4061 447
rect 4195 481 4319 487
rect 4195 447 4207 481
rect 4307 447 4319 481
rect 4195 441 4319 447
rect 4453 481 4577 487
rect 4453 447 4465 481
rect 4565 447 4577 481
rect 4453 441 4577 447
rect -4667 388 -4621 400
rect -4667 -388 -4661 388
rect -4627 -388 -4621 388
rect -4667 -400 -4621 -388
rect -4409 388 -4363 400
rect -4409 -388 -4403 388
rect -4369 -388 -4363 388
rect -4409 -400 -4363 -388
rect -4151 388 -4105 400
rect -4151 -388 -4145 388
rect -4111 -388 -4105 388
rect -4151 -400 -4105 -388
rect -3893 388 -3847 400
rect -3893 -388 -3887 388
rect -3853 -388 -3847 388
rect -3893 -400 -3847 -388
rect -3635 388 -3589 400
rect -3635 -388 -3629 388
rect -3595 -388 -3589 388
rect -3635 -400 -3589 -388
rect -3377 388 -3331 400
rect -3377 -388 -3371 388
rect -3337 -388 -3331 388
rect -3377 -400 -3331 -388
rect -3119 388 -3073 400
rect -3119 -388 -3113 388
rect -3079 -388 -3073 388
rect -3119 -400 -3073 -388
rect -2861 388 -2815 400
rect -2861 -388 -2855 388
rect -2821 -388 -2815 388
rect -2861 -400 -2815 -388
rect -2603 388 -2557 400
rect -2603 -388 -2597 388
rect -2563 -388 -2557 388
rect -2603 -400 -2557 -388
rect -2345 388 -2299 400
rect -2345 -388 -2339 388
rect -2305 -388 -2299 388
rect -2345 -400 -2299 -388
rect -2087 388 -2041 400
rect -2087 -388 -2081 388
rect -2047 -388 -2041 388
rect -2087 -400 -2041 -388
rect -1829 388 -1783 400
rect -1829 -388 -1823 388
rect -1789 -388 -1783 388
rect -1829 -400 -1783 -388
rect -1571 388 -1525 400
rect -1571 -388 -1565 388
rect -1531 -388 -1525 388
rect -1571 -400 -1525 -388
rect -1313 388 -1267 400
rect -1313 -388 -1307 388
rect -1273 -388 -1267 388
rect -1313 -400 -1267 -388
rect -1055 388 -1009 400
rect -1055 -388 -1049 388
rect -1015 -388 -1009 388
rect -1055 -400 -1009 -388
rect -797 388 -751 400
rect -797 -388 -791 388
rect -757 -388 -751 388
rect -797 -400 -751 -388
rect -539 388 -493 400
rect -539 -388 -533 388
rect -499 -388 -493 388
rect -539 -400 -493 -388
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect 493 388 539 400
rect 493 -388 499 388
rect 533 -388 539 388
rect 493 -400 539 -388
rect 751 388 797 400
rect 751 -388 757 388
rect 791 -388 797 388
rect 751 -400 797 -388
rect 1009 388 1055 400
rect 1009 -388 1015 388
rect 1049 -388 1055 388
rect 1009 -400 1055 -388
rect 1267 388 1313 400
rect 1267 -388 1273 388
rect 1307 -388 1313 388
rect 1267 -400 1313 -388
rect 1525 388 1571 400
rect 1525 -388 1531 388
rect 1565 -388 1571 388
rect 1525 -400 1571 -388
rect 1783 388 1829 400
rect 1783 -388 1789 388
rect 1823 -388 1829 388
rect 1783 -400 1829 -388
rect 2041 388 2087 400
rect 2041 -388 2047 388
rect 2081 -388 2087 388
rect 2041 -400 2087 -388
rect 2299 388 2345 400
rect 2299 -388 2305 388
rect 2339 -388 2345 388
rect 2299 -400 2345 -388
rect 2557 388 2603 400
rect 2557 -388 2563 388
rect 2597 -388 2603 388
rect 2557 -400 2603 -388
rect 2815 388 2861 400
rect 2815 -388 2821 388
rect 2855 -388 2861 388
rect 2815 -400 2861 -388
rect 3073 388 3119 400
rect 3073 -388 3079 388
rect 3113 -388 3119 388
rect 3073 -400 3119 -388
rect 3331 388 3377 400
rect 3331 -388 3337 388
rect 3371 -388 3377 388
rect 3331 -400 3377 -388
rect 3589 388 3635 400
rect 3589 -388 3595 388
rect 3629 -388 3635 388
rect 3589 -400 3635 -388
rect 3847 388 3893 400
rect 3847 -388 3853 388
rect 3887 -388 3893 388
rect 3847 -400 3893 -388
rect 4105 388 4151 400
rect 4105 -388 4111 388
rect 4145 -388 4151 388
rect 4105 -400 4151 -388
rect 4363 388 4409 400
rect 4363 -388 4369 388
rect 4403 -388 4409 388
rect 4363 -400 4409 -388
rect 4621 388 4667 400
rect 4621 -388 4627 388
rect 4661 -388 4667 388
rect 4621 -400 4667 -388
rect -4577 -447 -4453 -441
rect -4577 -481 -4565 -447
rect -4465 -481 -4453 -447
rect -4577 -487 -4453 -481
rect -4319 -447 -4195 -441
rect -4319 -481 -4307 -447
rect -4207 -481 -4195 -447
rect -4319 -487 -4195 -481
rect -4061 -447 -3937 -441
rect -4061 -481 -4049 -447
rect -3949 -481 -3937 -447
rect -4061 -487 -3937 -481
rect -3803 -447 -3679 -441
rect -3803 -481 -3791 -447
rect -3691 -481 -3679 -447
rect -3803 -487 -3679 -481
rect -3545 -447 -3421 -441
rect -3545 -481 -3533 -447
rect -3433 -481 -3421 -447
rect -3545 -487 -3421 -481
rect -3287 -447 -3163 -441
rect -3287 -481 -3275 -447
rect -3175 -481 -3163 -447
rect -3287 -487 -3163 -481
rect -3029 -447 -2905 -441
rect -3029 -481 -3017 -447
rect -2917 -481 -2905 -447
rect -3029 -487 -2905 -481
rect -2771 -447 -2647 -441
rect -2771 -481 -2759 -447
rect -2659 -481 -2647 -447
rect -2771 -487 -2647 -481
rect -2513 -447 -2389 -441
rect -2513 -481 -2501 -447
rect -2401 -481 -2389 -447
rect -2513 -487 -2389 -481
rect -2255 -447 -2131 -441
rect -2255 -481 -2243 -447
rect -2143 -481 -2131 -447
rect -2255 -487 -2131 -481
rect -1997 -447 -1873 -441
rect -1997 -481 -1985 -447
rect -1885 -481 -1873 -447
rect -1997 -487 -1873 -481
rect -1739 -447 -1615 -441
rect -1739 -481 -1727 -447
rect -1627 -481 -1615 -447
rect -1739 -487 -1615 -481
rect -1481 -447 -1357 -441
rect -1481 -481 -1469 -447
rect -1369 -481 -1357 -447
rect -1481 -487 -1357 -481
rect -1223 -447 -1099 -441
rect -1223 -481 -1211 -447
rect -1111 -481 -1099 -447
rect -1223 -487 -1099 -481
rect -965 -447 -841 -441
rect -965 -481 -953 -447
rect -853 -481 -841 -447
rect -965 -487 -841 -481
rect -707 -447 -583 -441
rect -707 -481 -695 -447
rect -595 -481 -583 -447
rect -707 -487 -583 -481
rect -449 -447 -325 -441
rect -449 -481 -437 -447
rect -337 -481 -325 -447
rect -449 -487 -325 -481
rect -191 -447 -67 -441
rect -191 -481 -179 -447
rect -79 -481 -67 -447
rect -191 -487 -67 -481
rect 67 -447 191 -441
rect 67 -481 79 -447
rect 179 -481 191 -447
rect 67 -487 191 -481
rect 325 -447 449 -441
rect 325 -481 337 -447
rect 437 -481 449 -447
rect 325 -487 449 -481
rect 583 -447 707 -441
rect 583 -481 595 -447
rect 695 -481 707 -447
rect 583 -487 707 -481
rect 841 -447 965 -441
rect 841 -481 853 -447
rect 953 -481 965 -447
rect 841 -487 965 -481
rect 1099 -447 1223 -441
rect 1099 -481 1111 -447
rect 1211 -481 1223 -447
rect 1099 -487 1223 -481
rect 1357 -447 1481 -441
rect 1357 -481 1369 -447
rect 1469 -481 1481 -447
rect 1357 -487 1481 -481
rect 1615 -447 1739 -441
rect 1615 -481 1627 -447
rect 1727 -481 1739 -447
rect 1615 -487 1739 -481
rect 1873 -447 1997 -441
rect 1873 -481 1885 -447
rect 1985 -481 1997 -447
rect 1873 -487 1997 -481
rect 2131 -447 2255 -441
rect 2131 -481 2143 -447
rect 2243 -481 2255 -447
rect 2131 -487 2255 -481
rect 2389 -447 2513 -441
rect 2389 -481 2401 -447
rect 2501 -481 2513 -447
rect 2389 -487 2513 -481
rect 2647 -447 2771 -441
rect 2647 -481 2659 -447
rect 2759 -481 2771 -447
rect 2647 -487 2771 -481
rect 2905 -447 3029 -441
rect 2905 -481 2917 -447
rect 3017 -481 3029 -447
rect 2905 -487 3029 -481
rect 3163 -447 3287 -441
rect 3163 -481 3175 -447
rect 3275 -481 3287 -447
rect 3163 -487 3287 -481
rect 3421 -447 3545 -441
rect 3421 -481 3433 -447
rect 3533 -481 3545 -447
rect 3421 -487 3545 -481
rect 3679 -447 3803 -441
rect 3679 -481 3691 -447
rect 3791 -481 3803 -447
rect 3679 -487 3803 -481
rect 3937 -447 4061 -441
rect 3937 -481 3949 -447
rect 4049 -481 4061 -447
rect 3937 -487 4061 -481
rect 4195 -447 4319 -441
rect 4195 -481 4207 -447
rect 4307 -481 4319 -447
rect 4195 -487 4319 -481
rect 4453 -447 4577 -441
rect 4453 -481 4465 -447
rect 4565 -481 4577 -447
rect 4453 -487 4577 -481
<< properties >>
string FIXED_BBOX -4778 -602 4778 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 36 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

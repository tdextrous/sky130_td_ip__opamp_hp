magic
tech sky130A
magscale 1 2
timestamp 1713234499
<< nwell >>
rect -1019 -1197 1019 1197
<< mvpmos >>
rect -761 -900 -661 900
rect -603 -900 -503 900
rect -445 -900 -345 900
rect -287 -900 -187 900
rect -129 -900 -29 900
rect 29 -900 129 900
rect 187 -900 287 900
rect 345 -900 445 900
rect 503 -900 603 900
rect 661 -900 761 900
<< mvpdiff >>
rect -819 888 -761 900
rect -819 -888 -807 888
rect -773 -888 -761 888
rect -819 -900 -761 -888
rect -661 888 -603 900
rect -661 -888 -649 888
rect -615 -888 -603 888
rect -661 -900 -603 -888
rect -503 888 -445 900
rect -503 -888 -491 888
rect -457 -888 -445 888
rect -503 -900 -445 -888
rect -345 888 -287 900
rect -345 -888 -333 888
rect -299 -888 -287 888
rect -345 -900 -287 -888
rect -187 888 -129 900
rect -187 -888 -175 888
rect -141 -888 -129 888
rect -187 -900 -129 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 129 888 187 900
rect 129 -888 141 888
rect 175 -888 187 888
rect 129 -900 187 -888
rect 287 888 345 900
rect 287 -888 299 888
rect 333 -888 345 888
rect 287 -900 345 -888
rect 445 888 503 900
rect 445 -888 457 888
rect 491 -888 503 888
rect 445 -900 503 -888
rect 603 888 661 900
rect 603 -888 615 888
rect 649 -888 661 888
rect 603 -900 661 -888
rect 761 888 819 900
rect 761 -888 773 888
rect 807 -888 819 888
rect 761 -900 819 -888
<< mvpdiffc >>
rect -807 -888 -773 888
rect -649 -888 -615 888
rect -491 -888 -457 888
rect -333 -888 -299 888
rect -175 -888 -141 888
rect -17 -888 17 888
rect 141 -888 175 888
rect 299 -888 333 888
rect 457 -888 491 888
rect 615 -888 649 888
rect 773 -888 807 888
<< mvnsubdiff >>
rect -953 1119 953 1131
rect -953 1085 -845 1119
rect 845 1085 953 1119
rect -953 1073 953 1085
rect -953 1023 -895 1073
rect -953 -1023 -941 1023
rect -907 -1023 -895 1023
rect 895 1023 953 1073
rect -953 -1073 -895 -1023
rect 895 -1023 907 1023
rect 941 -1023 953 1023
rect 895 -1073 953 -1023
rect -953 -1085 953 -1073
rect -953 -1119 -845 -1085
rect 845 -1119 953 -1085
rect -953 -1131 953 -1119
<< mvnsubdiffcont >>
rect -845 1085 845 1119
rect -941 -1023 -907 1023
rect 907 -1023 941 1023
rect -845 -1119 845 -1085
<< poly >>
rect -761 981 -661 997
rect -761 947 -745 981
rect -677 947 -661 981
rect -761 900 -661 947
rect -603 981 -503 997
rect -603 947 -587 981
rect -519 947 -503 981
rect -603 900 -503 947
rect -445 981 -345 997
rect -445 947 -429 981
rect -361 947 -345 981
rect -445 900 -345 947
rect -287 981 -187 997
rect -287 947 -271 981
rect -203 947 -187 981
rect -287 900 -187 947
rect -129 981 -29 997
rect -129 947 -113 981
rect -45 947 -29 981
rect -129 900 -29 947
rect 29 981 129 997
rect 29 947 45 981
rect 113 947 129 981
rect 29 900 129 947
rect 187 981 287 997
rect 187 947 203 981
rect 271 947 287 981
rect 187 900 287 947
rect 345 981 445 997
rect 345 947 361 981
rect 429 947 445 981
rect 345 900 445 947
rect 503 981 603 997
rect 503 947 519 981
rect 587 947 603 981
rect 503 900 603 947
rect 661 981 761 997
rect 661 947 677 981
rect 745 947 761 981
rect 661 900 761 947
rect -761 -947 -661 -900
rect -761 -981 -745 -947
rect -677 -981 -661 -947
rect -761 -997 -661 -981
rect -603 -947 -503 -900
rect -603 -981 -587 -947
rect -519 -981 -503 -947
rect -603 -997 -503 -981
rect -445 -947 -345 -900
rect -445 -981 -429 -947
rect -361 -981 -345 -947
rect -445 -997 -345 -981
rect -287 -947 -187 -900
rect -287 -981 -271 -947
rect -203 -981 -187 -947
rect -287 -997 -187 -981
rect -129 -947 -29 -900
rect -129 -981 -113 -947
rect -45 -981 -29 -947
rect -129 -997 -29 -981
rect 29 -947 129 -900
rect 29 -981 45 -947
rect 113 -981 129 -947
rect 29 -997 129 -981
rect 187 -947 287 -900
rect 187 -981 203 -947
rect 271 -981 287 -947
rect 187 -997 287 -981
rect 345 -947 445 -900
rect 345 -981 361 -947
rect 429 -981 445 -947
rect 345 -997 445 -981
rect 503 -947 603 -900
rect 503 -981 519 -947
rect 587 -981 603 -947
rect 503 -997 603 -981
rect 661 -947 761 -900
rect 661 -981 677 -947
rect 745 -981 761 -947
rect 661 -997 761 -981
<< polycont >>
rect -745 947 -677 981
rect -587 947 -519 981
rect -429 947 -361 981
rect -271 947 -203 981
rect -113 947 -45 981
rect 45 947 113 981
rect 203 947 271 981
rect 361 947 429 981
rect 519 947 587 981
rect 677 947 745 981
rect -745 -981 -677 -947
rect -587 -981 -519 -947
rect -429 -981 -361 -947
rect -271 -981 -203 -947
rect -113 -981 -45 -947
rect 45 -981 113 -947
rect 203 -981 271 -947
rect 361 -981 429 -947
rect 519 -981 587 -947
rect 677 -981 745 -947
<< locali >>
rect -941 1085 -845 1119
rect 845 1085 941 1119
rect -941 1023 -907 1085
rect 907 1023 941 1085
rect -761 947 -745 981
rect -677 947 -661 981
rect -603 947 -587 981
rect -519 947 -503 981
rect -445 947 -429 981
rect -361 947 -345 981
rect -287 947 -271 981
rect -203 947 -187 981
rect -129 947 -113 981
rect -45 947 -29 981
rect 29 947 45 981
rect 113 947 129 981
rect 187 947 203 981
rect 271 947 287 981
rect 345 947 361 981
rect 429 947 445 981
rect 503 947 519 981
rect 587 947 603 981
rect 661 947 677 981
rect 745 947 761 981
rect -807 888 -773 904
rect -807 -904 -773 -888
rect -649 888 -615 904
rect -649 -904 -615 -888
rect -491 888 -457 904
rect -491 -904 -457 -888
rect -333 888 -299 904
rect -333 -904 -299 -888
rect -175 888 -141 904
rect -175 -904 -141 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 141 888 175 904
rect 141 -904 175 -888
rect 299 888 333 904
rect 299 -904 333 -888
rect 457 888 491 904
rect 457 -904 491 -888
rect 615 888 649 904
rect 615 -904 649 -888
rect 773 888 807 904
rect 773 -904 807 -888
rect -761 -981 -745 -947
rect -677 -981 -661 -947
rect -603 -981 -587 -947
rect -519 -981 -503 -947
rect -445 -981 -429 -947
rect -361 -981 -345 -947
rect -287 -981 -271 -947
rect -203 -981 -187 -947
rect -129 -981 -113 -947
rect -45 -981 -29 -947
rect 29 -981 45 -947
rect 113 -981 129 -947
rect 187 -981 203 -947
rect 271 -981 287 -947
rect 345 -981 361 -947
rect 429 -981 445 -947
rect 503 -981 519 -947
rect 587 -981 603 -947
rect 661 -981 677 -947
rect 745 -981 761 -947
rect -941 -1085 -907 -1023
rect 907 -1085 941 -1023
rect -941 -1119 -845 -1085
rect 845 -1119 941 -1085
<< viali >>
rect -745 947 -677 981
rect -587 947 -519 981
rect -429 947 -361 981
rect -271 947 -203 981
rect -113 947 -45 981
rect 45 947 113 981
rect 203 947 271 981
rect 361 947 429 981
rect 519 947 587 981
rect 677 947 745 981
rect -807 -888 -773 888
rect -649 -888 -615 888
rect -491 -888 -457 888
rect -333 -888 -299 888
rect -175 -888 -141 888
rect -17 -888 17 888
rect 141 -888 175 888
rect 299 -888 333 888
rect 457 -888 491 888
rect 615 -888 649 888
rect 773 -888 807 888
rect -745 -981 -677 -947
rect -587 -981 -519 -947
rect -429 -981 -361 -947
rect -271 -981 -203 -947
rect -113 -981 -45 -947
rect 45 -981 113 -947
rect 203 -981 271 -947
rect 361 -981 429 -947
rect 519 -981 587 -947
rect 677 -981 745 -947
<< metal1 >>
rect -757 981 -665 987
rect -757 947 -745 981
rect -677 947 -665 981
rect -757 941 -665 947
rect -599 981 -507 987
rect -599 947 -587 981
rect -519 947 -507 981
rect -599 941 -507 947
rect -441 981 -349 987
rect -441 947 -429 981
rect -361 947 -349 981
rect -441 941 -349 947
rect -283 981 -191 987
rect -283 947 -271 981
rect -203 947 -191 981
rect -283 941 -191 947
rect -125 981 -33 987
rect -125 947 -113 981
rect -45 947 -33 981
rect -125 941 -33 947
rect 33 981 125 987
rect 33 947 45 981
rect 113 947 125 981
rect 33 941 125 947
rect 191 981 283 987
rect 191 947 203 981
rect 271 947 283 981
rect 191 941 283 947
rect 349 981 441 987
rect 349 947 361 981
rect 429 947 441 981
rect 349 941 441 947
rect 507 981 599 987
rect 507 947 519 981
rect 587 947 599 981
rect 507 941 599 947
rect 665 981 757 987
rect 665 947 677 981
rect 745 947 757 981
rect 665 941 757 947
rect -813 888 -767 900
rect -813 -888 -807 888
rect -773 -888 -767 888
rect -813 -900 -767 -888
rect -655 888 -609 900
rect -655 -888 -649 888
rect -615 -888 -609 888
rect -655 -900 -609 -888
rect -497 888 -451 900
rect -497 -888 -491 888
rect -457 -888 -451 888
rect -497 -900 -451 -888
rect -339 888 -293 900
rect -339 -888 -333 888
rect -299 -888 -293 888
rect -339 -900 -293 -888
rect -181 888 -135 900
rect -181 -888 -175 888
rect -141 -888 -135 888
rect -181 -900 -135 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 135 888 181 900
rect 135 -888 141 888
rect 175 -888 181 888
rect 135 -900 181 -888
rect 293 888 339 900
rect 293 -888 299 888
rect 333 -888 339 888
rect 293 -900 339 -888
rect 451 888 497 900
rect 451 -888 457 888
rect 491 -888 497 888
rect 451 -900 497 -888
rect 609 888 655 900
rect 609 -888 615 888
rect 649 -888 655 888
rect 609 -900 655 -888
rect 767 888 813 900
rect 767 -888 773 888
rect 807 -888 813 888
rect 767 -900 813 -888
rect -757 -947 -665 -941
rect -757 -981 -745 -947
rect -677 -981 -665 -947
rect -757 -987 -665 -981
rect -599 -947 -507 -941
rect -599 -981 -587 -947
rect -519 -981 -507 -947
rect -599 -987 -507 -981
rect -441 -947 -349 -941
rect -441 -981 -429 -947
rect -361 -981 -349 -947
rect -441 -987 -349 -981
rect -283 -947 -191 -941
rect -283 -981 -271 -947
rect -203 -981 -191 -947
rect -283 -987 -191 -981
rect -125 -947 -33 -941
rect -125 -981 -113 -947
rect -45 -981 -33 -947
rect -125 -987 -33 -981
rect 33 -947 125 -941
rect 33 -981 45 -947
rect 113 -981 125 -947
rect 33 -987 125 -981
rect 191 -947 283 -941
rect 191 -981 203 -947
rect 271 -981 283 -947
rect 191 -987 283 -981
rect 349 -947 441 -941
rect 349 -981 361 -947
rect 429 -981 441 -947
rect 349 -987 441 -981
rect 507 -947 599 -941
rect 507 -981 519 -947
rect 587 -981 599 -947
rect 507 -987 599 -981
rect 665 -947 757 -941
rect 665 -981 677 -947
rect 745 -981 757 -947
rect 665 -987 757 -981
<< properties >>
string FIXED_BBOX -924 -1102 924 1102
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

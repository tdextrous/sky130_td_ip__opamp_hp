magic
tech sky130A
magscale 1 2
timestamp 1713239177
<< pwell >>
rect -4585 -1258 4585 1258
<< mvnmos >>
rect -4357 -1000 -4157 1000
rect -4099 -1000 -3899 1000
rect -3841 -1000 -3641 1000
rect -3583 -1000 -3383 1000
rect -3325 -1000 -3125 1000
rect -3067 -1000 -2867 1000
rect -2809 -1000 -2609 1000
rect -2551 -1000 -2351 1000
rect -2293 -1000 -2093 1000
rect -2035 -1000 -1835 1000
rect -1777 -1000 -1577 1000
rect -1519 -1000 -1319 1000
rect -1261 -1000 -1061 1000
rect -1003 -1000 -803 1000
rect -745 -1000 -545 1000
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
rect 545 -1000 745 1000
rect 803 -1000 1003 1000
rect 1061 -1000 1261 1000
rect 1319 -1000 1519 1000
rect 1577 -1000 1777 1000
rect 1835 -1000 2035 1000
rect 2093 -1000 2293 1000
rect 2351 -1000 2551 1000
rect 2609 -1000 2809 1000
rect 2867 -1000 3067 1000
rect 3125 -1000 3325 1000
rect 3383 -1000 3583 1000
rect 3641 -1000 3841 1000
rect 3899 -1000 4099 1000
rect 4157 -1000 4357 1000
<< mvndiff >>
rect -4415 988 -4357 1000
rect -4415 -988 -4403 988
rect -4369 -988 -4357 988
rect -4415 -1000 -4357 -988
rect -4157 988 -4099 1000
rect -4157 -988 -4145 988
rect -4111 -988 -4099 988
rect -4157 -1000 -4099 -988
rect -3899 988 -3841 1000
rect -3899 -988 -3887 988
rect -3853 -988 -3841 988
rect -3899 -1000 -3841 -988
rect -3641 988 -3583 1000
rect -3641 -988 -3629 988
rect -3595 -988 -3583 988
rect -3641 -1000 -3583 -988
rect -3383 988 -3325 1000
rect -3383 -988 -3371 988
rect -3337 -988 -3325 988
rect -3383 -1000 -3325 -988
rect -3125 988 -3067 1000
rect -3125 -988 -3113 988
rect -3079 -988 -3067 988
rect -3125 -1000 -3067 -988
rect -2867 988 -2809 1000
rect -2867 -988 -2855 988
rect -2821 -988 -2809 988
rect -2867 -1000 -2809 -988
rect -2609 988 -2551 1000
rect -2609 -988 -2597 988
rect -2563 -988 -2551 988
rect -2609 -1000 -2551 -988
rect -2351 988 -2293 1000
rect -2351 -988 -2339 988
rect -2305 -988 -2293 988
rect -2351 -1000 -2293 -988
rect -2093 988 -2035 1000
rect -2093 -988 -2081 988
rect -2047 -988 -2035 988
rect -2093 -1000 -2035 -988
rect -1835 988 -1777 1000
rect -1835 -988 -1823 988
rect -1789 -988 -1777 988
rect -1835 -1000 -1777 -988
rect -1577 988 -1519 1000
rect -1577 -988 -1565 988
rect -1531 -988 -1519 988
rect -1577 -1000 -1519 -988
rect -1319 988 -1261 1000
rect -1319 -988 -1307 988
rect -1273 -988 -1261 988
rect -1319 -1000 -1261 -988
rect -1061 988 -1003 1000
rect -1061 -988 -1049 988
rect -1015 -988 -1003 988
rect -1061 -1000 -1003 -988
rect -803 988 -745 1000
rect -803 -988 -791 988
rect -757 -988 -745 988
rect -803 -1000 -745 -988
rect -545 988 -487 1000
rect -545 -988 -533 988
rect -499 -988 -487 988
rect -545 -1000 -487 -988
rect -287 988 -229 1000
rect -287 -988 -275 988
rect -241 -988 -229 988
rect -287 -1000 -229 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 229 988 287 1000
rect 229 -988 241 988
rect 275 -988 287 988
rect 229 -1000 287 -988
rect 487 988 545 1000
rect 487 -988 499 988
rect 533 -988 545 988
rect 487 -1000 545 -988
rect 745 988 803 1000
rect 745 -988 757 988
rect 791 -988 803 988
rect 745 -1000 803 -988
rect 1003 988 1061 1000
rect 1003 -988 1015 988
rect 1049 -988 1061 988
rect 1003 -1000 1061 -988
rect 1261 988 1319 1000
rect 1261 -988 1273 988
rect 1307 -988 1319 988
rect 1261 -1000 1319 -988
rect 1519 988 1577 1000
rect 1519 -988 1531 988
rect 1565 -988 1577 988
rect 1519 -1000 1577 -988
rect 1777 988 1835 1000
rect 1777 -988 1789 988
rect 1823 -988 1835 988
rect 1777 -1000 1835 -988
rect 2035 988 2093 1000
rect 2035 -988 2047 988
rect 2081 -988 2093 988
rect 2035 -1000 2093 -988
rect 2293 988 2351 1000
rect 2293 -988 2305 988
rect 2339 -988 2351 988
rect 2293 -1000 2351 -988
rect 2551 988 2609 1000
rect 2551 -988 2563 988
rect 2597 -988 2609 988
rect 2551 -1000 2609 -988
rect 2809 988 2867 1000
rect 2809 -988 2821 988
rect 2855 -988 2867 988
rect 2809 -1000 2867 -988
rect 3067 988 3125 1000
rect 3067 -988 3079 988
rect 3113 -988 3125 988
rect 3067 -1000 3125 -988
rect 3325 988 3383 1000
rect 3325 -988 3337 988
rect 3371 -988 3383 988
rect 3325 -1000 3383 -988
rect 3583 988 3641 1000
rect 3583 -988 3595 988
rect 3629 -988 3641 988
rect 3583 -1000 3641 -988
rect 3841 988 3899 1000
rect 3841 -988 3853 988
rect 3887 -988 3899 988
rect 3841 -1000 3899 -988
rect 4099 988 4157 1000
rect 4099 -988 4111 988
rect 4145 -988 4157 988
rect 4099 -1000 4157 -988
rect 4357 988 4415 1000
rect 4357 -988 4369 988
rect 4403 -988 4415 988
rect 4357 -1000 4415 -988
<< mvndiffc >>
rect -4403 -988 -4369 988
rect -4145 -988 -4111 988
rect -3887 -988 -3853 988
rect -3629 -988 -3595 988
rect -3371 -988 -3337 988
rect -3113 -988 -3079 988
rect -2855 -988 -2821 988
rect -2597 -988 -2563 988
rect -2339 -988 -2305 988
rect -2081 -988 -2047 988
rect -1823 -988 -1789 988
rect -1565 -988 -1531 988
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect 1531 -988 1565 988
rect 1789 -988 1823 988
rect 2047 -988 2081 988
rect 2305 -988 2339 988
rect 2563 -988 2597 988
rect 2821 -988 2855 988
rect 3079 -988 3113 988
rect 3337 -988 3371 988
rect 3595 -988 3629 988
rect 3853 -988 3887 988
rect 4111 -988 4145 988
rect 4369 -988 4403 988
<< mvpsubdiff >>
rect -4549 1210 4549 1222
rect -4549 1176 -4441 1210
rect 4441 1176 4549 1210
rect -4549 1164 4549 1176
rect -4549 1114 -4491 1164
rect -4549 -1114 -4537 1114
rect -4503 -1114 -4491 1114
rect 4491 1114 4549 1164
rect -4549 -1164 -4491 -1114
rect 4491 -1114 4503 1114
rect 4537 -1114 4549 1114
rect 4491 -1164 4549 -1114
rect -4549 -1176 4549 -1164
rect -4549 -1210 -4441 -1176
rect 4441 -1210 4549 -1176
rect -4549 -1222 4549 -1210
<< mvpsubdiffcont >>
rect -4441 1176 4441 1210
rect -4537 -1114 -4503 1114
rect 4503 -1114 4537 1114
rect -4441 -1210 4441 -1176
<< poly >>
rect -4357 1072 -4157 1088
rect -4357 1038 -4341 1072
rect -4173 1038 -4157 1072
rect -4357 1000 -4157 1038
rect -4099 1072 -3899 1088
rect -4099 1038 -4083 1072
rect -3915 1038 -3899 1072
rect -4099 1000 -3899 1038
rect -3841 1072 -3641 1088
rect -3841 1038 -3825 1072
rect -3657 1038 -3641 1072
rect -3841 1000 -3641 1038
rect -3583 1072 -3383 1088
rect -3583 1038 -3567 1072
rect -3399 1038 -3383 1072
rect -3583 1000 -3383 1038
rect -3325 1072 -3125 1088
rect -3325 1038 -3309 1072
rect -3141 1038 -3125 1072
rect -3325 1000 -3125 1038
rect -3067 1072 -2867 1088
rect -3067 1038 -3051 1072
rect -2883 1038 -2867 1072
rect -3067 1000 -2867 1038
rect -2809 1072 -2609 1088
rect -2809 1038 -2793 1072
rect -2625 1038 -2609 1072
rect -2809 1000 -2609 1038
rect -2551 1072 -2351 1088
rect -2551 1038 -2535 1072
rect -2367 1038 -2351 1072
rect -2551 1000 -2351 1038
rect -2293 1072 -2093 1088
rect -2293 1038 -2277 1072
rect -2109 1038 -2093 1072
rect -2293 1000 -2093 1038
rect -2035 1072 -1835 1088
rect -2035 1038 -2019 1072
rect -1851 1038 -1835 1072
rect -2035 1000 -1835 1038
rect -1777 1072 -1577 1088
rect -1777 1038 -1761 1072
rect -1593 1038 -1577 1072
rect -1777 1000 -1577 1038
rect -1519 1072 -1319 1088
rect -1519 1038 -1503 1072
rect -1335 1038 -1319 1072
rect -1519 1000 -1319 1038
rect -1261 1072 -1061 1088
rect -1261 1038 -1245 1072
rect -1077 1038 -1061 1072
rect -1261 1000 -1061 1038
rect -1003 1072 -803 1088
rect -1003 1038 -987 1072
rect -819 1038 -803 1072
rect -1003 1000 -803 1038
rect -745 1072 -545 1088
rect -745 1038 -729 1072
rect -561 1038 -545 1072
rect -745 1000 -545 1038
rect -487 1072 -287 1088
rect -487 1038 -471 1072
rect -303 1038 -287 1072
rect -487 1000 -287 1038
rect -229 1072 -29 1088
rect -229 1038 -213 1072
rect -45 1038 -29 1072
rect -229 1000 -29 1038
rect 29 1072 229 1088
rect 29 1038 45 1072
rect 213 1038 229 1072
rect 29 1000 229 1038
rect 287 1072 487 1088
rect 287 1038 303 1072
rect 471 1038 487 1072
rect 287 1000 487 1038
rect 545 1072 745 1088
rect 545 1038 561 1072
rect 729 1038 745 1072
rect 545 1000 745 1038
rect 803 1072 1003 1088
rect 803 1038 819 1072
rect 987 1038 1003 1072
rect 803 1000 1003 1038
rect 1061 1072 1261 1088
rect 1061 1038 1077 1072
rect 1245 1038 1261 1072
rect 1061 1000 1261 1038
rect 1319 1072 1519 1088
rect 1319 1038 1335 1072
rect 1503 1038 1519 1072
rect 1319 1000 1519 1038
rect 1577 1072 1777 1088
rect 1577 1038 1593 1072
rect 1761 1038 1777 1072
rect 1577 1000 1777 1038
rect 1835 1072 2035 1088
rect 1835 1038 1851 1072
rect 2019 1038 2035 1072
rect 1835 1000 2035 1038
rect 2093 1072 2293 1088
rect 2093 1038 2109 1072
rect 2277 1038 2293 1072
rect 2093 1000 2293 1038
rect 2351 1072 2551 1088
rect 2351 1038 2367 1072
rect 2535 1038 2551 1072
rect 2351 1000 2551 1038
rect 2609 1072 2809 1088
rect 2609 1038 2625 1072
rect 2793 1038 2809 1072
rect 2609 1000 2809 1038
rect 2867 1072 3067 1088
rect 2867 1038 2883 1072
rect 3051 1038 3067 1072
rect 2867 1000 3067 1038
rect 3125 1072 3325 1088
rect 3125 1038 3141 1072
rect 3309 1038 3325 1072
rect 3125 1000 3325 1038
rect 3383 1072 3583 1088
rect 3383 1038 3399 1072
rect 3567 1038 3583 1072
rect 3383 1000 3583 1038
rect 3641 1072 3841 1088
rect 3641 1038 3657 1072
rect 3825 1038 3841 1072
rect 3641 1000 3841 1038
rect 3899 1072 4099 1088
rect 3899 1038 3915 1072
rect 4083 1038 4099 1072
rect 3899 1000 4099 1038
rect 4157 1072 4357 1088
rect 4157 1038 4173 1072
rect 4341 1038 4357 1072
rect 4157 1000 4357 1038
rect -4357 -1038 -4157 -1000
rect -4357 -1072 -4341 -1038
rect -4173 -1072 -4157 -1038
rect -4357 -1088 -4157 -1072
rect -4099 -1038 -3899 -1000
rect -4099 -1072 -4083 -1038
rect -3915 -1072 -3899 -1038
rect -4099 -1088 -3899 -1072
rect -3841 -1038 -3641 -1000
rect -3841 -1072 -3825 -1038
rect -3657 -1072 -3641 -1038
rect -3841 -1088 -3641 -1072
rect -3583 -1038 -3383 -1000
rect -3583 -1072 -3567 -1038
rect -3399 -1072 -3383 -1038
rect -3583 -1088 -3383 -1072
rect -3325 -1038 -3125 -1000
rect -3325 -1072 -3309 -1038
rect -3141 -1072 -3125 -1038
rect -3325 -1088 -3125 -1072
rect -3067 -1038 -2867 -1000
rect -3067 -1072 -3051 -1038
rect -2883 -1072 -2867 -1038
rect -3067 -1088 -2867 -1072
rect -2809 -1038 -2609 -1000
rect -2809 -1072 -2793 -1038
rect -2625 -1072 -2609 -1038
rect -2809 -1088 -2609 -1072
rect -2551 -1038 -2351 -1000
rect -2551 -1072 -2535 -1038
rect -2367 -1072 -2351 -1038
rect -2551 -1088 -2351 -1072
rect -2293 -1038 -2093 -1000
rect -2293 -1072 -2277 -1038
rect -2109 -1072 -2093 -1038
rect -2293 -1088 -2093 -1072
rect -2035 -1038 -1835 -1000
rect -2035 -1072 -2019 -1038
rect -1851 -1072 -1835 -1038
rect -2035 -1088 -1835 -1072
rect -1777 -1038 -1577 -1000
rect -1777 -1072 -1761 -1038
rect -1593 -1072 -1577 -1038
rect -1777 -1088 -1577 -1072
rect -1519 -1038 -1319 -1000
rect -1519 -1072 -1503 -1038
rect -1335 -1072 -1319 -1038
rect -1519 -1088 -1319 -1072
rect -1261 -1038 -1061 -1000
rect -1261 -1072 -1245 -1038
rect -1077 -1072 -1061 -1038
rect -1261 -1088 -1061 -1072
rect -1003 -1038 -803 -1000
rect -1003 -1072 -987 -1038
rect -819 -1072 -803 -1038
rect -1003 -1088 -803 -1072
rect -745 -1038 -545 -1000
rect -745 -1072 -729 -1038
rect -561 -1072 -545 -1038
rect -745 -1088 -545 -1072
rect -487 -1038 -287 -1000
rect -487 -1072 -471 -1038
rect -303 -1072 -287 -1038
rect -487 -1088 -287 -1072
rect -229 -1038 -29 -1000
rect -229 -1072 -213 -1038
rect -45 -1072 -29 -1038
rect -229 -1088 -29 -1072
rect 29 -1038 229 -1000
rect 29 -1072 45 -1038
rect 213 -1072 229 -1038
rect 29 -1088 229 -1072
rect 287 -1038 487 -1000
rect 287 -1072 303 -1038
rect 471 -1072 487 -1038
rect 287 -1088 487 -1072
rect 545 -1038 745 -1000
rect 545 -1072 561 -1038
rect 729 -1072 745 -1038
rect 545 -1088 745 -1072
rect 803 -1038 1003 -1000
rect 803 -1072 819 -1038
rect 987 -1072 1003 -1038
rect 803 -1088 1003 -1072
rect 1061 -1038 1261 -1000
rect 1061 -1072 1077 -1038
rect 1245 -1072 1261 -1038
rect 1061 -1088 1261 -1072
rect 1319 -1038 1519 -1000
rect 1319 -1072 1335 -1038
rect 1503 -1072 1519 -1038
rect 1319 -1088 1519 -1072
rect 1577 -1038 1777 -1000
rect 1577 -1072 1593 -1038
rect 1761 -1072 1777 -1038
rect 1577 -1088 1777 -1072
rect 1835 -1038 2035 -1000
rect 1835 -1072 1851 -1038
rect 2019 -1072 2035 -1038
rect 1835 -1088 2035 -1072
rect 2093 -1038 2293 -1000
rect 2093 -1072 2109 -1038
rect 2277 -1072 2293 -1038
rect 2093 -1088 2293 -1072
rect 2351 -1038 2551 -1000
rect 2351 -1072 2367 -1038
rect 2535 -1072 2551 -1038
rect 2351 -1088 2551 -1072
rect 2609 -1038 2809 -1000
rect 2609 -1072 2625 -1038
rect 2793 -1072 2809 -1038
rect 2609 -1088 2809 -1072
rect 2867 -1038 3067 -1000
rect 2867 -1072 2883 -1038
rect 3051 -1072 3067 -1038
rect 2867 -1088 3067 -1072
rect 3125 -1038 3325 -1000
rect 3125 -1072 3141 -1038
rect 3309 -1072 3325 -1038
rect 3125 -1088 3325 -1072
rect 3383 -1038 3583 -1000
rect 3383 -1072 3399 -1038
rect 3567 -1072 3583 -1038
rect 3383 -1088 3583 -1072
rect 3641 -1038 3841 -1000
rect 3641 -1072 3657 -1038
rect 3825 -1072 3841 -1038
rect 3641 -1088 3841 -1072
rect 3899 -1038 4099 -1000
rect 3899 -1072 3915 -1038
rect 4083 -1072 4099 -1038
rect 3899 -1088 4099 -1072
rect 4157 -1038 4357 -1000
rect 4157 -1072 4173 -1038
rect 4341 -1072 4357 -1038
rect 4157 -1088 4357 -1072
<< polycont >>
rect -4341 1038 -4173 1072
rect -4083 1038 -3915 1072
rect -3825 1038 -3657 1072
rect -3567 1038 -3399 1072
rect -3309 1038 -3141 1072
rect -3051 1038 -2883 1072
rect -2793 1038 -2625 1072
rect -2535 1038 -2367 1072
rect -2277 1038 -2109 1072
rect -2019 1038 -1851 1072
rect -1761 1038 -1593 1072
rect -1503 1038 -1335 1072
rect -1245 1038 -1077 1072
rect -987 1038 -819 1072
rect -729 1038 -561 1072
rect -471 1038 -303 1072
rect -213 1038 -45 1072
rect 45 1038 213 1072
rect 303 1038 471 1072
rect 561 1038 729 1072
rect 819 1038 987 1072
rect 1077 1038 1245 1072
rect 1335 1038 1503 1072
rect 1593 1038 1761 1072
rect 1851 1038 2019 1072
rect 2109 1038 2277 1072
rect 2367 1038 2535 1072
rect 2625 1038 2793 1072
rect 2883 1038 3051 1072
rect 3141 1038 3309 1072
rect 3399 1038 3567 1072
rect 3657 1038 3825 1072
rect 3915 1038 4083 1072
rect 4173 1038 4341 1072
rect -4341 -1072 -4173 -1038
rect -4083 -1072 -3915 -1038
rect -3825 -1072 -3657 -1038
rect -3567 -1072 -3399 -1038
rect -3309 -1072 -3141 -1038
rect -3051 -1072 -2883 -1038
rect -2793 -1072 -2625 -1038
rect -2535 -1072 -2367 -1038
rect -2277 -1072 -2109 -1038
rect -2019 -1072 -1851 -1038
rect -1761 -1072 -1593 -1038
rect -1503 -1072 -1335 -1038
rect -1245 -1072 -1077 -1038
rect -987 -1072 -819 -1038
rect -729 -1072 -561 -1038
rect -471 -1072 -303 -1038
rect -213 -1072 -45 -1038
rect 45 -1072 213 -1038
rect 303 -1072 471 -1038
rect 561 -1072 729 -1038
rect 819 -1072 987 -1038
rect 1077 -1072 1245 -1038
rect 1335 -1072 1503 -1038
rect 1593 -1072 1761 -1038
rect 1851 -1072 2019 -1038
rect 2109 -1072 2277 -1038
rect 2367 -1072 2535 -1038
rect 2625 -1072 2793 -1038
rect 2883 -1072 3051 -1038
rect 3141 -1072 3309 -1038
rect 3399 -1072 3567 -1038
rect 3657 -1072 3825 -1038
rect 3915 -1072 4083 -1038
rect 4173 -1072 4341 -1038
<< locali >>
rect -4537 1176 -4441 1210
rect 4441 1176 4537 1210
rect -4537 1114 -4503 1176
rect 4503 1114 4537 1176
rect -4357 1038 -4341 1072
rect -4173 1038 -4157 1072
rect -4099 1038 -4083 1072
rect -3915 1038 -3899 1072
rect -3841 1038 -3825 1072
rect -3657 1038 -3641 1072
rect -3583 1038 -3567 1072
rect -3399 1038 -3383 1072
rect -3325 1038 -3309 1072
rect -3141 1038 -3125 1072
rect -3067 1038 -3051 1072
rect -2883 1038 -2867 1072
rect -2809 1038 -2793 1072
rect -2625 1038 -2609 1072
rect -2551 1038 -2535 1072
rect -2367 1038 -2351 1072
rect -2293 1038 -2277 1072
rect -2109 1038 -2093 1072
rect -2035 1038 -2019 1072
rect -1851 1038 -1835 1072
rect -1777 1038 -1761 1072
rect -1593 1038 -1577 1072
rect -1519 1038 -1503 1072
rect -1335 1038 -1319 1072
rect -1261 1038 -1245 1072
rect -1077 1038 -1061 1072
rect -1003 1038 -987 1072
rect -819 1038 -803 1072
rect -745 1038 -729 1072
rect -561 1038 -545 1072
rect -487 1038 -471 1072
rect -303 1038 -287 1072
rect -229 1038 -213 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 213 1038 229 1072
rect 287 1038 303 1072
rect 471 1038 487 1072
rect 545 1038 561 1072
rect 729 1038 745 1072
rect 803 1038 819 1072
rect 987 1038 1003 1072
rect 1061 1038 1077 1072
rect 1245 1038 1261 1072
rect 1319 1038 1335 1072
rect 1503 1038 1519 1072
rect 1577 1038 1593 1072
rect 1761 1038 1777 1072
rect 1835 1038 1851 1072
rect 2019 1038 2035 1072
rect 2093 1038 2109 1072
rect 2277 1038 2293 1072
rect 2351 1038 2367 1072
rect 2535 1038 2551 1072
rect 2609 1038 2625 1072
rect 2793 1038 2809 1072
rect 2867 1038 2883 1072
rect 3051 1038 3067 1072
rect 3125 1038 3141 1072
rect 3309 1038 3325 1072
rect 3383 1038 3399 1072
rect 3567 1038 3583 1072
rect 3641 1038 3657 1072
rect 3825 1038 3841 1072
rect 3899 1038 3915 1072
rect 4083 1038 4099 1072
rect 4157 1038 4173 1072
rect 4341 1038 4357 1072
rect -4403 988 -4369 1004
rect -4403 -1004 -4369 -988
rect -4145 988 -4111 1004
rect -4145 -1004 -4111 -988
rect -3887 988 -3853 1004
rect -3887 -1004 -3853 -988
rect -3629 988 -3595 1004
rect -3629 -1004 -3595 -988
rect -3371 988 -3337 1004
rect -3371 -1004 -3337 -988
rect -3113 988 -3079 1004
rect -3113 -1004 -3079 -988
rect -2855 988 -2821 1004
rect -2855 -1004 -2821 -988
rect -2597 988 -2563 1004
rect -2597 -1004 -2563 -988
rect -2339 988 -2305 1004
rect -2339 -1004 -2305 -988
rect -2081 988 -2047 1004
rect -2081 -1004 -2047 -988
rect -1823 988 -1789 1004
rect -1823 -1004 -1789 -988
rect -1565 988 -1531 1004
rect -1565 -1004 -1531 -988
rect -1307 988 -1273 1004
rect -1307 -1004 -1273 -988
rect -1049 988 -1015 1004
rect -1049 -1004 -1015 -988
rect -791 988 -757 1004
rect -791 -1004 -757 -988
rect -533 988 -499 1004
rect -533 -1004 -499 -988
rect -275 988 -241 1004
rect -275 -1004 -241 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 241 988 275 1004
rect 241 -1004 275 -988
rect 499 988 533 1004
rect 499 -1004 533 -988
rect 757 988 791 1004
rect 757 -1004 791 -988
rect 1015 988 1049 1004
rect 1015 -1004 1049 -988
rect 1273 988 1307 1004
rect 1273 -1004 1307 -988
rect 1531 988 1565 1004
rect 1531 -1004 1565 -988
rect 1789 988 1823 1004
rect 1789 -1004 1823 -988
rect 2047 988 2081 1004
rect 2047 -1004 2081 -988
rect 2305 988 2339 1004
rect 2305 -1004 2339 -988
rect 2563 988 2597 1004
rect 2563 -1004 2597 -988
rect 2821 988 2855 1004
rect 2821 -1004 2855 -988
rect 3079 988 3113 1004
rect 3079 -1004 3113 -988
rect 3337 988 3371 1004
rect 3337 -1004 3371 -988
rect 3595 988 3629 1004
rect 3595 -1004 3629 -988
rect 3853 988 3887 1004
rect 3853 -1004 3887 -988
rect 4111 988 4145 1004
rect 4111 -1004 4145 -988
rect 4369 988 4403 1004
rect 4369 -1004 4403 -988
rect -4357 -1072 -4341 -1038
rect -4173 -1072 -4157 -1038
rect -4099 -1072 -4083 -1038
rect -3915 -1072 -3899 -1038
rect -3841 -1072 -3825 -1038
rect -3657 -1072 -3641 -1038
rect -3583 -1072 -3567 -1038
rect -3399 -1072 -3383 -1038
rect -3325 -1072 -3309 -1038
rect -3141 -1072 -3125 -1038
rect -3067 -1072 -3051 -1038
rect -2883 -1072 -2867 -1038
rect -2809 -1072 -2793 -1038
rect -2625 -1072 -2609 -1038
rect -2551 -1072 -2535 -1038
rect -2367 -1072 -2351 -1038
rect -2293 -1072 -2277 -1038
rect -2109 -1072 -2093 -1038
rect -2035 -1072 -2019 -1038
rect -1851 -1072 -1835 -1038
rect -1777 -1072 -1761 -1038
rect -1593 -1072 -1577 -1038
rect -1519 -1072 -1503 -1038
rect -1335 -1072 -1319 -1038
rect -1261 -1072 -1245 -1038
rect -1077 -1072 -1061 -1038
rect -1003 -1072 -987 -1038
rect -819 -1072 -803 -1038
rect -745 -1072 -729 -1038
rect -561 -1072 -545 -1038
rect -487 -1072 -471 -1038
rect -303 -1072 -287 -1038
rect -229 -1072 -213 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 213 -1072 229 -1038
rect 287 -1072 303 -1038
rect 471 -1072 487 -1038
rect 545 -1072 561 -1038
rect 729 -1072 745 -1038
rect 803 -1072 819 -1038
rect 987 -1072 1003 -1038
rect 1061 -1072 1077 -1038
rect 1245 -1072 1261 -1038
rect 1319 -1072 1335 -1038
rect 1503 -1072 1519 -1038
rect 1577 -1072 1593 -1038
rect 1761 -1072 1777 -1038
rect 1835 -1072 1851 -1038
rect 2019 -1072 2035 -1038
rect 2093 -1072 2109 -1038
rect 2277 -1072 2293 -1038
rect 2351 -1072 2367 -1038
rect 2535 -1072 2551 -1038
rect 2609 -1072 2625 -1038
rect 2793 -1072 2809 -1038
rect 2867 -1072 2883 -1038
rect 3051 -1072 3067 -1038
rect 3125 -1072 3141 -1038
rect 3309 -1072 3325 -1038
rect 3383 -1072 3399 -1038
rect 3567 -1072 3583 -1038
rect 3641 -1072 3657 -1038
rect 3825 -1072 3841 -1038
rect 3899 -1072 3915 -1038
rect 4083 -1072 4099 -1038
rect 4157 -1072 4173 -1038
rect 4341 -1072 4357 -1038
rect -4537 -1176 -4503 -1114
rect 4503 -1176 4537 -1114
rect -4537 -1210 -4441 -1176
rect 4441 -1210 4537 -1176
<< viali >>
rect -4341 1038 -4173 1072
rect -4083 1038 -3915 1072
rect -3825 1038 -3657 1072
rect -3567 1038 -3399 1072
rect -3309 1038 -3141 1072
rect -3051 1038 -2883 1072
rect -2793 1038 -2625 1072
rect -2535 1038 -2367 1072
rect -2277 1038 -2109 1072
rect -2019 1038 -1851 1072
rect -1761 1038 -1593 1072
rect -1503 1038 -1335 1072
rect -1245 1038 -1077 1072
rect -987 1038 -819 1072
rect -729 1038 -561 1072
rect -471 1038 -303 1072
rect -213 1038 -45 1072
rect 45 1038 213 1072
rect 303 1038 471 1072
rect 561 1038 729 1072
rect 819 1038 987 1072
rect 1077 1038 1245 1072
rect 1335 1038 1503 1072
rect 1593 1038 1761 1072
rect 1851 1038 2019 1072
rect 2109 1038 2277 1072
rect 2367 1038 2535 1072
rect 2625 1038 2793 1072
rect 2883 1038 3051 1072
rect 3141 1038 3309 1072
rect 3399 1038 3567 1072
rect 3657 1038 3825 1072
rect 3915 1038 4083 1072
rect 4173 1038 4341 1072
rect -4403 -988 -4369 988
rect -4145 -988 -4111 988
rect -3887 -988 -3853 988
rect -3629 -988 -3595 988
rect -3371 -988 -3337 988
rect -3113 -988 -3079 988
rect -2855 -988 -2821 988
rect -2597 -988 -2563 988
rect -2339 -988 -2305 988
rect -2081 -988 -2047 988
rect -1823 -988 -1789 988
rect -1565 -988 -1531 988
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect 1531 -988 1565 988
rect 1789 -988 1823 988
rect 2047 -988 2081 988
rect 2305 -988 2339 988
rect 2563 -988 2597 988
rect 2821 -988 2855 988
rect 3079 -988 3113 988
rect 3337 -988 3371 988
rect 3595 -988 3629 988
rect 3853 -988 3887 988
rect 4111 -988 4145 988
rect 4369 -988 4403 988
rect -4341 -1072 -4173 -1038
rect -4083 -1072 -3915 -1038
rect -3825 -1072 -3657 -1038
rect -3567 -1072 -3399 -1038
rect -3309 -1072 -3141 -1038
rect -3051 -1072 -2883 -1038
rect -2793 -1072 -2625 -1038
rect -2535 -1072 -2367 -1038
rect -2277 -1072 -2109 -1038
rect -2019 -1072 -1851 -1038
rect -1761 -1072 -1593 -1038
rect -1503 -1072 -1335 -1038
rect -1245 -1072 -1077 -1038
rect -987 -1072 -819 -1038
rect -729 -1072 -561 -1038
rect -471 -1072 -303 -1038
rect -213 -1072 -45 -1038
rect 45 -1072 213 -1038
rect 303 -1072 471 -1038
rect 561 -1072 729 -1038
rect 819 -1072 987 -1038
rect 1077 -1072 1245 -1038
rect 1335 -1072 1503 -1038
rect 1593 -1072 1761 -1038
rect 1851 -1072 2019 -1038
rect 2109 -1072 2277 -1038
rect 2367 -1072 2535 -1038
rect 2625 -1072 2793 -1038
rect 2883 -1072 3051 -1038
rect 3141 -1072 3309 -1038
rect 3399 -1072 3567 -1038
rect 3657 -1072 3825 -1038
rect 3915 -1072 4083 -1038
rect 4173 -1072 4341 -1038
<< metal1 >>
rect -4353 1072 -4161 1078
rect -4353 1038 -4341 1072
rect -4173 1038 -4161 1072
rect -4353 1032 -4161 1038
rect -4095 1072 -3903 1078
rect -4095 1038 -4083 1072
rect -3915 1038 -3903 1072
rect -4095 1032 -3903 1038
rect -3837 1072 -3645 1078
rect -3837 1038 -3825 1072
rect -3657 1038 -3645 1072
rect -3837 1032 -3645 1038
rect -3579 1072 -3387 1078
rect -3579 1038 -3567 1072
rect -3399 1038 -3387 1072
rect -3579 1032 -3387 1038
rect -3321 1072 -3129 1078
rect -3321 1038 -3309 1072
rect -3141 1038 -3129 1072
rect -3321 1032 -3129 1038
rect -3063 1072 -2871 1078
rect -3063 1038 -3051 1072
rect -2883 1038 -2871 1072
rect -3063 1032 -2871 1038
rect -2805 1072 -2613 1078
rect -2805 1038 -2793 1072
rect -2625 1038 -2613 1072
rect -2805 1032 -2613 1038
rect -2547 1072 -2355 1078
rect -2547 1038 -2535 1072
rect -2367 1038 -2355 1072
rect -2547 1032 -2355 1038
rect -2289 1072 -2097 1078
rect -2289 1038 -2277 1072
rect -2109 1038 -2097 1072
rect -2289 1032 -2097 1038
rect -2031 1072 -1839 1078
rect -2031 1038 -2019 1072
rect -1851 1038 -1839 1072
rect -2031 1032 -1839 1038
rect -1773 1072 -1581 1078
rect -1773 1038 -1761 1072
rect -1593 1038 -1581 1072
rect -1773 1032 -1581 1038
rect -1515 1072 -1323 1078
rect -1515 1038 -1503 1072
rect -1335 1038 -1323 1072
rect -1515 1032 -1323 1038
rect -1257 1072 -1065 1078
rect -1257 1038 -1245 1072
rect -1077 1038 -1065 1072
rect -1257 1032 -1065 1038
rect -999 1072 -807 1078
rect -999 1038 -987 1072
rect -819 1038 -807 1072
rect -999 1032 -807 1038
rect -741 1072 -549 1078
rect -741 1038 -729 1072
rect -561 1038 -549 1072
rect -741 1032 -549 1038
rect -483 1072 -291 1078
rect -483 1038 -471 1072
rect -303 1038 -291 1072
rect -483 1032 -291 1038
rect -225 1072 -33 1078
rect -225 1038 -213 1072
rect -45 1038 -33 1072
rect -225 1032 -33 1038
rect 33 1072 225 1078
rect 33 1038 45 1072
rect 213 1038 225 1072
rect 33 1032 225 1038
rect 291 1072 483 1078
rect 291 1038 303 1072
rect 471 1038 483 1072
rect 291 1032 483 1038
rect 549 1072 741 1078
rect 549 1038 561 1072
rect 729 1038 741 1072
rect 549 1032 741 1038
rect 807 1072 999 1078
rect 807 1038 819 1072
rect 987 1038 999 1072
rect 807 1032 999 1038
rect 1065 1072 1257 1078
rect 1065 1038 1077 1072
rect 1245 1038 1257 1072
rect 1065 1032 1257 1038
rect 1323 1072 1515 1078
rect 1323 1038 1335 1072
rect 1503 1038 1515 1072
rect 1323 1032 1515 1038
rect 1581 1072 1773 1078
rect 1581 1038 1593 1072
rect 1761 1038 1773 1072
rect 1581 1032 1773 1038
rect 1839 1072 2031 1078
rect 1839 1038 1851 1072
rect 2019 1038 2031 1072
rect 1839 1032 2031 1038
rect 2097 1072 2289 1078
rect 2097 1038 2109 1072
rect 2277 1038 2289 1072
rect 2097 1032 2289 1038
rect 2355 1072 2547 1078
rect 2355 1038 2367 1072
rect 2535 1038 2547 1072
rect 2355 1032 2547 1038
rect 2613 1072 2805 1078
rect 2613 1038 2625 1072
rect 2793 1038 2805 1072
rect 2613 1032 2805 1038
rect 2871 1072 3063 1078
rect 2871 1038 2883 1072
rect 3051 1038 3063 1072
rect 2871 1032 3063 1038
rect 3129 1072 3321 1078
rect 3129 1038 3141 1072
rect 3309 1038 3321 1072
rect 3129 1032 3321 1038
rect 3387 1072 3579 1078
rect 3387 1038 3399 1072
rect 3567 1038 3579 1072
rect 3387 1032 3579 1038
rect 3645 1072 3837 1078
rect 3645 1038 3657 1072
rect 3825 1038 3837 1072
rect 3645 1032 3837 1038
rect 3903 1072 4095 1078
rect 3903 1038 3915 1072
rect 4083 1038 4095 1072
rect 3903 1032 4095 1038
rect 4161 1072 4353 1078
rect 4161 1038 4173 1072
rect 4341 1038 4353 1072
rect 4161 1032 4353 1038
rect -4409 988 -4363 1000
rect -4409 -988 -4403 988
rect -4369 -988 -4363 988
rect -4409 -1000 -4363 -988
rect -4151 988 -4105 1000
rect -4151 -988 -4145 988
rect -4111 -988 -4105 988
rect -4151 -1000 -4105 -988
rect -3893 988 -3847 1000
rect -3893 -988 -3887 988
rect -3853 -988 -3847 988
rect -3893 -1000 -3847 -988
rect -3635 988 -3589 1000
rect -3635 -988 -3629 988
rect -3595 -988 -3589 988
rect -3635 -1000 -3589 -988
rect -3377 988 -3331 1000
rect -3377 -988 -3371 988
rect -3337 -988 -3331 988
rect -3377 -1000 -3331 -988
rect -3119 988 -3073 1000
rect -3119 -988 -3113 988
rect -3079 -988 -3073 988
rect -3119 -1000 -3073 -988
rect -2861 988 -2815 1000
rect -2861 -988 -2855 988
rect -2821 -988 -2815 988
rect -2861 -1000 -2815 -988
rect -2603 988 -2557 1000
rect -2603 -988 -2597 988
rect -2563 -988 -2557 988
rect -2603 -1000 -2557 -988
rect -2345 988 -2299 1000
rect -2345 -988 -2339 988
rect -2305 -988 -2299 988
rect -2345 -1000 -2299 -988
rect -2087 988 -2041 1000
rect -2087 -988 -2081 988
rect -2047 -988 -2041 988
rect -2087 -1000 -2041 -988
rect -1829 988 -1783 1000
rect -1829 -988 -1823 988
rect -1789 -988 -1783 988
rect -1829 -1000 -1783 -988
rect -1571 988 -1525 1000
rect -1571 -988 -1565 988
rect -1531 -988 -1525 988
rect -1571 -1000 -1525 -988
rect -1313 988 -1267 1000
rect -1313 -988 -1307 988
rect -1273 -988 -1267 988
rect -1313 -1000 -1267 -988
rect -1055 988 -1009 1000
rect -1055 -988 -1049 988
rect -1015 -988 -1009 988
rect -1055 -1000 -1009 -988
rect -797 988 -751 1000
rect -797 -988 -791 988
rect -757 -988 -751 988
rect -797 -1000 -751 -988
rect -539 988 -493 1000
rect -539 -988 -533 988
rect -499 -988 -493 988
rect -539 -1000 -493 -988
rect -281 988 -235 1000
rect -281 -988 -275 988
rect -241 -988 -235 988
rect -281 -1000 -235 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 235 988 281 1000
rect 235 -988 241 988
rect 275 -988 281 988
rect 235 -1000 281 -988
rect 493 988 539 1000
rect 493 -988 499 988
rect 533 -988 539 988
rect 493 -1000 539 -988
rect 751 988 797 1000
rect 751 -988 757 988
rect 791 -988 797 988
rect 751 -1000 797 -988
rect 1009 988 1055 1000
rect 1009 -988 1015 988
rect 1049 -988 1055 988
rect 1009 -1000 1055 -988
rect 1267 988 1313 1000
rect 1267 -988 1273 988
rect 1307 -988 1313 988
rect 1267 -1000 1313 -988
rect 1525 988 1571 1000
rect 1525 -988 1531 988
rect 1565 -988 1571 988
rect 1525 -1000 1571 -988
rect 1783 988 1829 1000
rect 1783 -988 1789 988
rect 1823 -988 1829 988
rect 1783 -1000 1829 -988
rect 2041 988 2087 1000
rect 2041 -988 2047 988
rect 2081 -988 2087 988
rect 2041 -1000 2087 -988
rect 2299 988 2345 1000
rect 2299 -988 2305 988
rect 2339 -988 2345 988
rect 2299 -1000 2345 -988
rect 2557 988 2603 1000
rect 2557 -988 2563 988
rect 2597 -988 2603 988
rect 2557 -1000 2603 -988
rect 2815 988 2861 1000
rect 2815 -988 2821 988
rect 2855 -988 2861 988
rect 2815 -1000 2861 -988
rect 3073 988 3119 1000
rect 3073 -988 3079 988
rect 3113 -988 3119 988
rect 3073 -1000 3119 -988
rect 3331 988 3377 1000
rect 3331 -988 3337 988
rect 3371 -988 3377 988
rect 3331 -1000 3377 -988
rect 3589 988 3635 1000
rect 3589 -988 3595 988
rect 3629 -988 3635 988
rect 3589 -1000 3635 -988
rect 3847 988 3893 1000
rect 3847 -988 3853 988
rect 3887 -988 3893 988
rect 3847 -1000 3893 -988
rect 4105 988 4151 1000
rect 4105 -988 4111 988
rect 4145 -988 4151 988
rect 4105 -1000 4151 -988
rect 4363 988 4409 1000
rect 4363 -988 4369 988
rect 4403 -988 4409 988
rect 4363 -1000 4409 -988
rect -4353 -1038 -4161 -1032
rect -4353 -1072 -4341 -1038
rect -4173 -1072 -4161 -1038
rect -4353 -1078 -4161 -1072
rect -4095 -1038 -3903 -1032
rect -4095 -1072 -4083 -1038
rect -3915 -1072 -3903 -1038
rect -4095 -1078 -3903 -1072
rect -3837 -1038 -3645 -1032
rect -3837 -1072 -3825 -1038
rect -3657 -1072 -3645 -1038
rect -3837 -1078 -3645 -1072
rect -3579 -1038 -3387 -1032
rect -3579 -1072 -3567 -1038
rect -3399 -1072 -3387 -1038
rect -3579 -1078 -3387 -1072
rect -3321 -1038 -3129 -1032
rect -3321 -1072 -3309 -1038
rect -3141 -1072 -3129 -1038
rect -3321 -1078 -3129 -1072
rect -3063 -1038 -2871 -1032
rect -3063 -1072 -3051 -1038
rect -2883 -1072 -2871 -1038
rect -3063 -1078 -2871 -1072
rect -2805 -1038 -2613 -1032
rect -2805 -1072 -2793 -1038
rect -2625 -1072 -2613 -1038
rect -2805 -1078 -2613 -1072
rect -2547 -1038 -2355 -1032
rect -2547 -1072 -2535 -1038
rect -2367 -1072 -2355 -1038
rect -2547 -1078 -2355 -1072
rect -2289 -1038 -2097 -1032
rect -2289 -1072 -2277 -1038
rect -2109 -1072 -2097 -1038
rect -2289 -1078 -2097 -1072
rect -2031 -1038 -1839 -1032
rect -2031 -1072 -2019 -1038
rect -1851 -1072 -1839 -1038
rect -2031 -1078 -1839 -1072
rect -1773 -1038 -1581 -1032
rect -1773 -1072 -1761 -1038
rect -1593 -1072 -1581 -1038
rect -1773 -1078 -1581 -1072
rect -1515 -1038 -1323 -1032
rect -1515 -1072 -1503 -1038
rect -1335 -1072 -1323 -1038
rect -1515 -1078 -1323 -1072
rect -1257 -1038 -1065 -1032
rect -1257 -1072 -1245 -1038
rect -1077 -1072 -1065 -1038
rect -1257 -1078 -1065 -1072
rect -999 -1038 -807 -1032
rect -999 -1072 -987 -1038
rect -819 -1072 -807 -1038
rect -999 -1078 -807 -1072
rect -741 -1038 -549 -1032
rect -741 -1072 -729 -1038
rect -561 -1072 -549 -1038
rect -741 -1078 -549 -1072
rect -483 -1038 -291 -1032
rect -483 -1072 -471 -1038
rect -303 -1072 -291 -1038
rect -483 -1078 -291 -1072
rect -225 -1038 -33 -1032
rect -225 -1072 -213 -1038
rect -45 -1072 -33 -1038
rect -225 -1078 -33 -1072
rect 33 -1038 225 -1032
rect 33 -1072 45 -1038
rect 213 -1072 225 -1038
rect 33 -1078 225 -1072
rect 291 -1038 483 -1032
rect 291 -1072 303 -1038
rect 471 -1072 483 -1038
rect 291 -1078 483 -1072
rect 549 -1038 741 -1032
rect 549 -1072 561 -1038
rect 729 -1072 741 -1038
rect 549 -1078 741 -1072
rect 807 -1038 999 -1032
rect 807 -1072 819 -1038
rect 987 -1072 999 -1038
rect 807 -1078 999 -1072
rect 1065 -1038 1257 -1032
rect 1065 -1072 1077 -1038
rect 1245 -1072 1257 -1038
rect 1065 -1078 1257 -1072
rect 1323 -1038 1515 -1032
rect 1323 -1072 1335 -1038
rect 1503 -1072 1515 -1038
rect 1323 -1078 1515 -1072
rect 1581 -1038 1773 -1032
rect 1581 -1072 1593 -1038
rect 1761 -1072 1773 -1038
rect 1581 -1078 1773 -1072
rect 1839 -1038 2031 -1032
rect 1839 -1072 1851 -1038
rect 2019 -1072 2031 -1038
rect 1839 -1078 2031 -1072
rect 2097 -1038 2289 -1032
rect 2097 -1072 2109 -1038
rect 2277 -1072 2289 -1038
rect 2097 -1078 2289 -1072
rect 2355 -1038 2547 -1032
rect 2355 -1072 2367 -1038
rect 2535 -1072 2547 -1038
rect 2355 -1078 2547 -1072
rect 2613 -1038 2805 -1032
rect 2613 -1072 2625 -1038
rect 2793 -1072 2805 -1038
rect 2613 -1078 2805 -1072
rect 2871 -1038 3063 -1032
rect 2871 -1072 2883 -1038
rect 3051 -1072 3063 -1038
rect 2871 -1078 3063 -1072
rect 3129 -1038 3321 -1032
rect 3129 -1072 3141 -1038
rect 3309 -1072 3321 -1038
rect 3129 -1078 3321 -1072
rect 3387 -1038 3579 -1032
rect 3387 -1072 3399 -1038
rect 3567 -1072 3579 -1038
rect 3387 -1078 3579 -1072
rect 3645 -1038 3837 -1032
rect 3645 -1072 3657 -1038
rect 3825 -1072 3837 -1038
rect 3645 -1078 3837 -1072
rect 3903 -1038 4095 -1032
rect 3903 -1072 3915 -1038
rect 4083 -1072 4095 -1038
rect 3903 -1078 4095 -1072
rect 4161 -1038 4353 -1032
rect 4161 -1072 4173 -1038
rect 4341 -1072 4353 -1038
rect 4161 -1078 4353 -1072
<< properties >>
string FIXED_BBOX -4520 -1193 4520 1193
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10 l 1 m 1 nf 34 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

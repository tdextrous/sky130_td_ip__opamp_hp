magic
tech sky130A
magscale 1 2
timestamp 1713233265
<< pwell >>
rect -673 -1158 673 1158
<< mvnmos >>
rect -445 -900 -345 900
rect -287 -900 -187 900
rect -129 -900 -29 900
rect 29 -900 129 900
rect 187 -900 287 900
rect 345 -900 445 900
<< mvndiff >>
rect -503 888 -445 900
rect -503 -888 -491 888
rect -457 -888 -445 888
rect -503 -900 -445 -888
rect -345 888 -287 900
rect -345 -888 -333 888
rect -299 -888 -287 888
rect -345 -900 -287 -888
rect -187 888 -129 900
rect -187 -888 -175 888
rect -141 -888 -129 888
rect -187 -900 -129 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 129 888 187 900
rect 129 -888 141 888
rect 175 -888 187 888
rect 129 -900 187 -888
rect 287 888 345 900
rect 287 -888 299 888
rect 333 -888 345 888
rect 287 -900 345 -888
rect 445 888 503 900
rect 445 -888 457 888
rect 491 -888 503 888
rect 445 -900 503 -888
<< mvndiffc >>
rect -491 -888 -457 888
rect -333 -888 -299 888
rect -175 -888 -141 888
rect -17 -888 17 888
rect 141 -888 175 888
rect 299 -888 333 888
rect 457 -888 491 888
<< mvpsubdiff >>
rect -637 1110 637 1122
rect -637 1076 -529 1110
rect 529 1076 637 1110
rect -637 1064 637 1076
rect -637 1014 -579 1064
rect -637 -1014 -625 1014
rect -591 -1014 -579 1014
rect 579 1014 637 1064
rect -637 -1064 -579 -1014
rect 579 -1014 591 1014
rect 625 -1014 637 1014
rect 579 -1064 637 -1014
rect -637 -1076 637 -1064
rect -637 -1110 -529 -1076
rect 529 -1110 637 -1076
rect -637 -1122 637 -1110
<< mvpsubdiffcont >>
rect -529 1076 529 1110
rect -625 -1014 -591 1014
rect 591 -1014 625 1014
rect -529 -1110 529 -1076
<< poly >>
rect -445 972 -345 988
rect -445 938 -429 972
rect -361 938 -345 972
rect -445 900 -345 938
rect -287 972 -187 988
rect -287 938 -271 972
rect -203 938 -187 972
rect -287 900 -187 938
rect -129 972 -29 988
rect -129 938 -113 972
rect -45 938 -29 972
rect -129 900 -29 938
rect 29 972 129 988
rect 29 938 45 972
rect 113 938 129 972
rect 29 900 129 938
rect 187 972 287 988
rect 187 938 203 972
rect 271 938 287 972
rect 187 900 287 938
rect 345 972 445 988
rect 345 938 361 972
rect 429 938 445 972
rect 345 900 445 938
rect -445 -938 -345 -900
rect -445 -972 -429 -938
rect -361 -972 -345 -938
rect -445 -988 -345 -972
rect -287 -938 -187 -900
rect -287 -972 -271 -938
rect -203 -972 -187 -938
rect -287 -988 -187 -972
rect -129 -938 -29 -900
rect -129 -972 -113 -938
rect -45 -972 -29 -938
rect -129 -988 -29 -972
rect 29 -938 129 -900
rect 29 -972 45 -938
rect 113 -972 129 -938
rect 29 -988 129 -972
rect 187 -938 287 -900
rect 187 -972 203 -938
rect 271 -972 287 -938
rect 187 -988 287 -972
rect 345 -938 445 -900
rect 345 -972 361 -938
rect 429 -972 445 -938
rect 345 -988 445 -972
<< polycont >>
rect -429 938 -361 972
rect -271 938 -203 972
rect -113 938 -45 972
rect 45 938 113 972
rect 203 938 271 972
rect 361 938 429 972
rect -429 -972 -361 -938
rect -271 -972 -203 -938
rect -113 -972 -45 -938
rect 45 -972 113 -938
rect 203 -972 271 -938
rect 361 -972 429 -938
<< locali >>
rect -625 1076 -529 1110
rect 529 1076 625 1110
rect -625 1014 -591 1076
rect 591 1014 625 1076
rect -445 938 -429 972
rect -361 938 -345 972
rect -287 938 -271 972
rect -203 938 -187 972
rect -129 938 -113 972
rect -45 938 -29 972
rect 29 938 45 972
rect 113 938 129 972
rect 187 938 203 972
rect 271 938 287 972
rect 345 938 361 972
rect 429 938 445 972
rect -491 888 -457 904
rect -491 -904 -457 -888
rect -333 888 -299 904
rect -333 -904 -299 -888
rect -175 888 -141 904
rect -175 -904 -141 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 141 888 175 904
rect 141 -904 175 -888
rect 299 888 333 904
rect 299 -904 333 -888
rect 457 888 491 904
rect 457 -904 491 -888
rect -445 -972 -429 -938
rect -361 -972 -345 -938
rect -287 -972 -271 -938
rect -203 -972 -187 -938
rect -129 -972 -113 -938
rect -45 -972 -29 -938
rect 29 -972 45 -938
rect 113 -972 129 -938
rect 187 -972 203 -938
rect 271 -972 287 -938
rect 345 -972 361 -938
rect 429 -972 445 -938
rect -625 -1076 -591 -1014
rect 591 -1076 625 -1014
rect -625 -1110 -529 -1076
rect 529 -1110 625 -1076
<< viali >>
rect -429 938 -361 972
rect -271 938 -203 972
rect -113 938 -45 972
rect 45 938 113 972
rect 203 938 271 972
rect 361 938 429 972
rect -491 -888 -457 888
rect -333 -888 -299 888
rect -175 -888 -141 888
rect -17 -888 17 888
rect 141 -888 175 888
rect 299 -888 333 888
rect 457 -888 491 888
rect -429 -972 -361 -938
rect -271 -972 -203 -938
rect -113 -972 -45 -938
rect 45 -972 113 -938
rect 203 -972 271 -938
rect 361 -972 429 -938
<< metal1 >>
rect -441 972 -349 978
rect -441 938 -429 972
rect -361 938 -349 972
rect -441 932 -349 938
rect -283 972 -191 978
rect -283 938 -271 972
rect -203 938 -191 972
rect -283 932 -191 938
rect -125 972 -33 978
rect -125 938 -113 972
rect -45 938 -33 972
rect -125 932 -33 938
rect 33 972 125 978
rect 33 938 45 972
rect 113 938 125 972
rect 33 932 125 938
rect 191 972 283 978
rect 191 938 203 972
rect 271 938 283 972
rect 191 932 283 938
rect 349 972 441 978
rect 349 938 361 972
rect 429 938 441 972
rect 349 932 441 938
rect -497 888 -451 900
rect -497 -888 -491 888
rect -457 -888 -451 888
rect -497 -900 -451 -888
rect -339 888 -293 900
rect -339 -888 -333 888
rect -299 -888 -293 888
rect -339 -900 -293 -888
rect -181 888 -135 900
rect -181 -888 -175 888
rect -141 -888 -135 888
rect -181 -900 -135 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 135 888 181 900
rect 135 -888 141 888
rect 175 -888 181 888
rect 135 -900 181 -888
rect 293 888 339 900
rect 293 -888 299 888
rect 333 -888 339 888
rect 293 -900 339 -888
rect 451 888 497 900
rect 451 -888 457 888
rect 491 -888 497 888
rect 451 -900 497 -888
rect -441 -938 -349 -932
rect -441 -972 -429 -938
rect -361 -972 -349 -938
rect -441 -978 -349 -972
rect -283 -938 -191 -932
rect -283 -972 -271 -938
rect -203 -972 -191 -938
rect -283 -978 -191 -972
rect -125 -938 -33 -932
rect -125 -972 -113 -938
rect -45 -972 -33 -938
rect -125 -978 -33 -972
rect 33 -938 125 -932
rect 33 -972 45 -938
rect 113 -972 125 -938
rect 33 -978 125 -972
rect 191 -938 283 -932
rect 191 -972 203 -938
rect 271 -972 283 -938
rect 191 -978 283 -972
rect 349 -938 441 -932
rect 349 -972 361 -938
rect 429 -972 441 -938
rect 349 -978 441 -972
<< properties >>
string FIXED_BBOX -608 -1093 608 1093
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 9 l 0.5 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

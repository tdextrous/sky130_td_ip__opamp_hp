magic
tech sky130A
magscale 1 2
timestamp 1713234499
<< pwell >>
rect -831 -708 831 708
<< mvnmos >>
rect -603 -450 -503 450
rect -445 -450 -345 450
rect -287 -450 -187 450
rect -129 -450 -29 450
rect 29 -450 129 450
rect 187 -450 287 450
rect 345 -450 445 450
rect 503 -450 603 450
<< mvndiff >>
rect -661 438 -603 450
rect -661 -438 -649 438
rect -615 -438 -603 438
rect -661 -450 -603 -438
rect -503 438 -445 450
rect -503 -438 -491 438
rect -457 -438 -445 438
rect -503 -450 -445 -438
rect -345 438 -287 450
rect -345 -438 -333 438
rect -299 -438 -287 438
rect -345 -450 -287 -438
rect -187 438 -129 450
rect -187 -438 -175 438
rect -141 -438 -129 438
rect -187 -450 -129 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 129 438 187 450
rect 129 -438 141 438
rect 175 -438 187 438
rect 129 -450 187 -438
rect 287 438 345 450
rect 287 -438 299 438
rect 333 -438 345 438
rect 287 -450 345 -438
rect 445 438 503 450
rect 445 -438 457 438
rect 491 -438 503 438
rect 445 -450 503 -438
rect 603 438 661 450
rect 603 -438 615 438
rect 649 -438 661 438
rect 603 -450 661 -438
<< mvndiffc >>
rect -649 -438 -615 438
rect -491 -438 -457 438
rect -333 -438 -299 438
rect -175 -438 -141 438
rect -17 -438 17 438
rect 141 -438 175 438
rect 299 -438 333 438
rect 457 -438 491 438
rect 615 -438 649 438
<< mvpsubdiff >>
rect -795 660 795 672
rect -795 626 -687 660
rect 687 626 795 660
rect -795 614 795 626
rect -795 564 -737 614
rect -795 -564 -783 564
rect -749 -564 -737 564
rect 737 564 795 614
rect -795 -614 -737 -564
rect 737 -564 749 564
rect 783 -564 795 564
rect 737 -614 795 -564
rect -795 -626 795 -614
rect -795 -660 -687 -626
rect 687 -660 795 -626
rect -795 -672 795 -660
<< mvpsubdiffcont >>
rect -687 626 687 660
rect -783 -564 -749 564
rect 749 -564 783 564
rect -687 -660 687 -626
<< poly >>
rect -603 522 -503 538
rect -603 488 -587 522
rect -519 488 -503 522
rect -603 450 -503 488
rect -445 522 -345 538
rect -445 488 -429 522
rect -361 488 -345 522
rect -445 450 -345 488
rect -287 522 -187 538
rect -287 488 -271 522
rect -203 488 -187 522
rect -287 450 -187 488
rect -129 522 -29 538
rect -129 488 -113 522
rect -45 488 -29 522
rect -129 450 -29 488
rect 29 522 129 538
rect 29 488 45 522
rect 113 488 129 522
rect 29 450 129 488
rect 187 522 287 538
rect 187 488 203 522
rect 271 488 287 522
rect 187 450 287 488
rect 345 522 445 538
rect 345 488 361 522
rect 429 488 445 522
rect 345 450 445 488
rect 503 522 603 538
rect 503 488 519 522
rect 587 488 603 522
rect 503 450 603 488
rect -603 -488 -503 -450
rect -603 -522 -587 -488
rect -519 -522 -503 -488
rect -603 -538 -503 -522
rect -445 -488 -345 -450
rect -445 -522 -429 -488
rect -361 -522 -345 -488
rect -445 -538 -345 -522
rect -287 -488 -187 -450
rect -287 -522 -271 -488
rect -203 -522 -187 -488
rect -287 -538 -187 -522
rect -129 -488 -29 -450
rect -129 -522 -113 -488
rect -45 -522 -29 -488
rect -129 -538 -29 -522
rect 29 -488 129 -450
rect 29 -522 45 -488
rect 113 -522 129 -488
rect 29 -538 129 -522
rect 187 -488 287 -450
rect 187 -522 203 -488
rect 271 -522 287 -488
rect 187 -538 287 -522
rect 345 -488 445 -450
rect 345 -522 361 -488
rect 429 -522 445 -488
rect 345 -538 445 -522
rect 503 -488 603 -450
rect 503 -522 519 -488
rect 587 -522 603 -488
rect 503 -538 603 -522
<< polycont >>
rect -587 488 -519 522
rect -429 488 -361 522
rect -271 488 -203 522
rect -113 488 -45 522
rect 45 488 113 522
rect 203 488 271 522
rect 361 488 429 522
rect 519 488 587 522
rect -587 -522 -519 -488
rect -429 -522 -361 -488
rect -271 -522 -203 -488
rect -113 -522 -45 -488
rect 45 -522 113 -488
rect 203 -522 271 -488
rect 361 -522 429 -488
rect 519 -522 587 -488
<< locali >>
rect -783 626 -687 660
rect 687 626 783 660
rect -783 564 -749 626
rect 749 564 783 626
rect -603 488 -587 522
rect -519 488 -503 522
rect -445 488 -429 522
rect -361 488 -345 522
rect -287 488 -271 522
rect -203 488 -187 522
rect -129 488 -113 522
rect -45 488 -29 522
rect 29 488 45 522
rect 113 488 129 522
rect 187 488 203 522
rect 271 488 287 522
rect 345 488 361 522
rect 429 488 445 522
rect 503 488 519 522
rect 587 488 603 522
rect -649 438 -615 454
rect -649 -454 -615 -438
rect -491 438 -457 454
rect -491 -454 -457 -438
rect -333 438 -299 454
rect -333 -454 -299 -438
rect -175 438 -141 454
rect -175 -454 -141 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 141 438 175 454
rect 141 -454 175 -438
rect 299 438 333 454
rect 299 -454 333 -438
rect 457 438 491 454
rect 457 -454 491 -438
rect 615 438 649 454
rect 615 -454 649 -438
rect -603 -522 -587 -488
rect -519 -522 -503 -488
rect -445 -522 -429 -488
rect -361 -522 -345 -488
rect -287 -522 -271 -488
rect -203 -522 -187 -488
rect -129 -522 -113 -488
rect -45 -522 -29 -488
rect 29 -522 45 -488
rect 113 -522 129 -488
rect 187 -522 203 -488
rect 271 -522 287 -488
rect 345 -522 361 -488
rect 429 -522 445 -488
rect 503 -522 519 -488
rect 587 -522 603 -488
rect -783 -626 -749 -564
rect 749 -626 783 -564
rect -783 -660 -687 -626
rect 687 -660 783 -626
<< viali >>
rect -587 488 -519 522
rect -429 488 -361 522
rect -271 488 -203 522
rect -113 488 -45 522
rect 45 488 113 522
rect 203 488 271 522
rect 361 488 429 522
rect 519 488 587 522
rect -649 -438 -615 438
rect -491 -438 -457 438
rect -333 -438 -299 438
rect -175 -438 -141 438
rect -17 -438 17 438
rect 141 -438 175 438
rect 299 -438 333 438
rect 457 -438 491 438
rect 615 -438 649 438
rect -587 -522 -519 -488
rect -429 -522 -361 -488
rect -271 -522 -203 -488
rect -113 -522 -45 -488
rect 45 -522 113 -488
rect 203 -522 271 -488
rect 361 -522 429 -488
rect 519 -522 587 -488
<< metal1 >>
rect -599 522 -507 528
rect -599 488 -587 522
rect -519 488 -507 522
rect -599 482 -507 488
rect -441 522 -349 528
rect -441 488 -429 522
rect -361 488 -349 522
rect -441 482 -349 488
rect -283 522 -191 528
rect -283 488 -271 522
rect -203 488 -191 522
rect -283 482 -191 488
rect -125 522 -33 528
rect -125 488 -113 522
rect -45 488 -33 522
rect -125 482 -33 488
rect 33 522 125 528
rect 33 488 45 522
rect 113 488 125 522
rect 33 482 125 488
rect 191 522 283 528
rect 191 488 203 522
rect 271 488 283 522
rect 191 482 283 488
rect 349 522 441 528
rect 349 488 361 522
rect 429 488 441 522
rect 349 482 441 488
rect 507 522 599 528
rect 507 488 519 522
rect 587 488 599 522
rect 507 482 599 488
rect -655 438 -609 450
rect -655 -438 -649 438
rect -615 -438 -609 438
rect -655 -450 -609 -438
rect -497 438 -451 450
rect -497 -438 -491 438
rect -457 -438 -451 438
rect -497 -450 -451 -438
rect -339 438 -293 450
rect -339 -438 -333 438
rect -299 -438 -293 438
rect -339 -450 -293 -438
rect -181 438 -135 450
rect -181 -438 -175 438
rect -141 -438 -135 438
rect -181 -450 -135 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 135 438 181 450
rect 135 -438 141 438
rect 175 -438 181 438
rect 135 -450 181 -438
rect 293 438 339 450
rect 293 -438 299 438
rect 333 -438 339 438
rect 293 -450 339 -438
rect 451 438 497 450
rect 451 -438 457 438
rect 491 -438 497 438
rect 451 -450 497 -438
rect 609 438 655 450
rect 609 -438 615 438
rect 649 -438 655 438
rect 609 -450 655 -438
rect -599 -488 -507 -482
rect -599 -522 -587 -488
rect -519 -522 -507 -488
rect -599 -528 -507 -522
rect -441 -488 -349 -482
rect -441 -522 -429 -488
rect -361 -522 -349 -488
rect -441 -528 -349 -522
rect -283 -488 -191 -482
rect -283 -522 -271 -488
rect -203 -522 -191 -488
rect -283 -528 -191 -522
rect -125 -488 -33 -482
rect -125 -522 -113 -488
rect -45 -522 -33 -488
rect -125 -528 -33 -522
rect 33 -488 125 -482
rect 33 -522 45 -488
rect 113 -522 125 -488
rect 33 -528 125 -522
rect 191 -488 283 -482
rect 191 -522 203 -488
rect 271 -522 283 -488
rect 191 -528 283 -522
rect 349 -488 441 -482
rect 349 -522 361 -488
rect 429 -522 441 -488
rect 349 -528 441 -522
rect 507 -488 599 -482
rect 507 -522 519 -488
rect 587 -522 599 -488
rect 507 -528 599 -522
<< properties >>
string FIXED_BBOX -766 -643 766 643
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713485303
<< dnwell >>
rect -7206 -6487 50963 15919
<< nwell >>
rect -7286 15713 51043 15999
rect -7286 -6281 -7000 15713
rect -3830 3045 33507 13150
rect 50757 -6281 51043 15713
rect -7286 -6567 51043 -6281
<< psubdiff >>
rect -7255 16137 -7231 16199
rect 51034 16137 51058 16199
rect -7705 15968 -7592 15992
rect -7705 -6464 -7592 -6440
rect 51264 15918 51327 15942
rect 51264 -6694 51327 -6670
rect -7710 -6929 -7686 -6803
rect 51106 -6929 51130 -6803
<< nsubdiff >>
rect -7249 15942 51006 15962
rect -7249 15908 -7169 15942
rect 50926 15908 51006 15942
rect -7249 15888 51006 15908
rect -7249 15882 -7175 15888
rect -7249 -6450 -7229 15882
rect -7195 -6450 -7175 15882
rect 50932 15882 51006 15888
rect -3776 13038 -3716 13072
rect 33385 13038 33445 13072
rect -3776 13012 -3742 13038
rect -3776 3122 -3742 3148
rect 33411 13012 33445 13038
rect 33411 3122 33445 3148
rect -3776 3088 -3716 3122
rect 33385 3088 33445 3122
rect -7249 -6456 -7175 -6450
rect 50932 -6450 50952 15882
rect 50986 -6450 51006 15882
rect 50932 -6456 51006 -6450
rect -7249 -6476 51006 -6456
rect -7249 -6510 -7169 -6476
rect 50926 -6510 51006 -6476
rect -7249 -6530 51006 -6510
<< mvpsubdiff >>
rect -6426 2651 -6346 2675
rect 33295 2502 33427 2526
rect 33295 -4887 33427 -4863
rect -6426 -5148 -6346 -5124
rect -6230 -5589 -6206 -5410
rect 33230 -5589 33254 -5410
<< psubdiffcont >>
rect -7231 16137 51034 16199
rect -7705 -6440 -7592 15968
rect 51264 -6670 51327 15918
rect -7686 -6929 51106 -6803
<< nsubdiffcont >>
rect -7169 15908 50926 15942
rect -7229 -6450 -7195 15882
rect -3716 13038 33385 13072
rect -3776 3148 -3742 13012
rect 33411 3148 33445 13012
rect -3716 3088 33385 3122
rect 50952 -6450 50986 15882
rect -7169 -6510 50926 -6476
<< mvpsubdiffcont >>
rect -6426 -5124 -6346 2651
rect 33295 -4863 33427 2502
rect -6206 -5589 33230 -5410
<< locali >>
rect -7704 16198 -7592 16206
rect 51032 16199 51330 16202
rect -7247 16198 -7231 16199
rect -7704 16140 -7231 16198
rect -7704 15984 -7592 16140
rect -7247 16137 -7231 16140
rect 51034 16138 51330 16199
rect 51034 16137 51050 16138
rect -7705 15968 -7592 15984
rect -9952 5157 -8224 5161
rect -9952 4985 -9948 5157
rect -9418 4985 -8224 5157
rect -9952 4979 -8224 4985
rect -9444 4411 -9316 4811
rect -8622 4417 -8496 4811
rect -9468 3781 -9324 3981
rect -8636 3777 -8494 3977
rect -9966 3626 -8238 3627
rect -9966 3623 -7705 3626
rect -9966 3449 -9960 3623
rect -9336 3449 -7705 3623
rect -9966 3445 -7705 3449
rect -8304 3444 -7705 3445
rect -7724 -6440 -7705 -6344
rect -7724 -6456 -7592 -6440
rect -7229 15908 -7169 15942
rect 50926 15908 50986 15942
rect -7229 15882 -7195 15908
rect -3777 15882 50986 15908
rect -3777 15092 50952 15882
rect -3777 14843 -3384 15092
rect -3768 14434 -3384 14843
rect 33104 14434 50952 15092
rect -3768 14155 50952 14434
rect -3768 13075 33378 14155
rect -3768 13072 33445 13075
rect -3776 13038 -3716 13072
rect 33385 13038 33445 13072
rect -3776 13012 33445 13038
rect -3742 12894 33411 13012
rect -3742 12882 12812 12894
rect -3742 12735 12006 12882
rect -3742 9129 -2366 12735
rect -1900 9129 -1850 12735
rect -1384 9129 -1334 12735
rect -868 9129 -818 12735
rect -654 12570 -510 12622
rect -352 9129 -302 12735
rect 164 9130 214 12735
rect 680 9129 730 12735
rect 1196 9129 1246 12735
rect 1712 12617 12006 12735
rect 1712 12609 9413 12617
rect 1712 10415 3354 12609
rect 3820 10415 3870 12609
rect 4336 10416 4386 12609
rect 4852 10415 4902 12609
rect 5368 10415 5418 12609
rect 5884 10415 5934 12609
rect 6400 10415 6450 12609
rect 6916 10415 6966 12609
rect 7432 10415 7482 12609
rect 7948 10415 7998 12609
rect 8464 12416 9413 12609
rect 9580 12456 9656 12617
rect 11002 12448 11080 12617
rect 8464 10608 9576 12416
rect 11250 12414 12006 12617
rect 11092 11682 12006 12414
rect 12414 11686 12812 12882
rect 13248 12760 33411 12894
rect 13248 12751 23704 12760
rect 13248 12566 13529 12751
rect 13725 12593 13951 12751
rect 13248 12151 13698 12566
rect 13248 11968 13529 12151
rect 13903 12120 13951 12593
rect 13729 11968 13951 12120
rect 14419 11968 14467 12751
rect 14935 11968 14983 12751
rect 15451 11968 15499 12751
rect 15967 11968 16015 12751
rect 16483 12594 16707 12751
rect 16890 12731 23704 12751
rect 16890 12730 22792 12731
rect 16483 12121 16531 12594
rect 16890 12564 17746 12730
rect 17926 12583 18061 12730
rect 18699 12582 19095 12730
rect 21281 12582 21415 12730
rect 16734 12549 17746 12564
rect 16734 12146 17891 12549
rect 16890 12137 17891 12146
rect 16483 11968 16709 12121
rect 16890 11968 17746 12137
rect 18872 12105 18923 12582
rect 21599 12548 22792 12730
rect 23267 12591 23704 12731
rect 23872 12621 24007 12760
rect 23267 12548 23836 12591
rect 21452 12137 22792 12548
rect 13248 11954 17746 11968
rect 17926 11954 18061 12102
rect 18701 11954 19094 12105
rect 21282 11954 21416 12103
rect 21599 11954 22792 12137
rect 13248 11757 22792 11954
rect 23137 11937 23836 12548
rect 23267 11778 23836 11937
rect 23267 11757 23704 11778
rect 13248 11686 23704 11757
rect 12414 11682 23704 11686
rect 11092 11608 23704 11682
rect 23872 11608 24008 11744
rect 24046 11608 24092 12760
rect 24562 11611 24608 12760
rect 24900 12609 25301 12760
rect 25077 11780 25126 12609
rect 24903 11611 25299 11780
rect 25594 11611 25640 12760
rect 26110 11611 26156 12760
rect 26626 11611 26672 12760
rect 27142 11611 27188 12760
rect 27658 11611 27704 12760
rect 28174 11611 28220 12760
rect 28690 11611 28736 12760
rect 29206 11611 29252 12760
rect 29722 11611 29768 12760
rect 30238 11611 30284 12760
rect 30754 11611 30800 12760
rect 31270 11611 31316 12760
rect 31609 12616 32011 12760
rect 31782 11775 31838 12616
rect 31612 11611 32010 11775
rect 32302 11611 32348 12760
rect 32818 11611 32864 12760
rect 32900 12623 33038 12760
rect 33203 12592 33411 12760
rect 33072 11772 33411 12592
rect 24425 11610 32864 11611
rect 32901 11610 33039 11744
rect 33203 11610 33411 11772
rect 24425 11608 33411 11610
rect 11092 11333 33411 11608
rect 8464 10415 9413 10608
rect 11092 10606 12186 11333
rect 1712 10414 9413 10415
rect 9582 10414 9656 10570
rect 11002 10414 11080 10568
rect 11250 10414 12186 10606
rect 1712 9654 12186 10414
rect 1712 9646 8933 9654
rect 1712 9129 3260 9646
rect 4402 9488 4812 9646
rect -3742 8232 3260 9129
rect -3742 8054 -1400 8232
rect -1006 8230 3260 8232
rect -3742 5930 -1276 8054
rect -3742 4758 -3292 5930
rect -2010 4758 -1276 5930
rect -3742 4748 -1276 4758
rect -3742 4744 -2362 4748
rect -3742 4702 -2992 4744
rect -2936 4742 -2362 4744
rect -2936 4702 -2680 4742
rect -3742 4700 -2680 4702
rect -2624 4706 -2362 4742
rect -2306 4706 -1276 4748
rect -2624 4700 -1276 4706
rect -3742 4536 -1276 4700
rect -3742 4530 -2110 4536
rect -3742 3342 -3570 4530
rect -3164 4346 -2110 4530
rect -3164 4334 -1978 4346
rect -3298 3544 -1978 4334
rect -1704 3624 -1276 4536
rect -3298 3536 -2110 3544
rect -3164 3348 -2110 3536
rect -1704 3446 -1400 3624
rect -1006 3446 -504 8230
rect -1704 3444 -504 3446
rect -220 3444 46 8230
rect 318 8228 3260 8230
rect 318 3444 884 8228
rect -1704 3442 884 3444
rect 1162 7456 3260 8228
rect 4576 7624 4644 9488
rect 9052 8532 12186 9654
rect 12482 8532 12528 11333
rect 12996 8532 13046 11333
rect 13084 11180 13100 11214
rect 13200 11180 13216 11214
rect 13342 11180 13358 11214
rect 13458 11180 13474 11214
rect 13262 11121 13296 11137
rect 13262 8729 13296 8745
rect 13084 8652 13100 8686
rect 13200 8652 13216 8686
rect 13342 8652 13358 8686
rect 13458 8652 13474 8686
rect 13512 8532 13562 11333
rect 14028 8532 14078 11333
rect 14116 11180 14132 11214
rect 14232 11180 14248 11214
rect 14374 11180 14390 11214
rect 14490 11180 14506 11214
rect 14294 11121 14328 11137
rect 14294 8729 14328 8745
rect 14116 8652 14132 8686
rect 14232 8652 14248 8686
rect 14374 8652 14390 8686
rect 14490 8652 14506 8686
rect 14544 8532 14594 11333
rect 14632 11180 14648 11214
rect 14748 11180 14764 11214
rect 14890 11180 14906 11214
rect 15006 11180 15022 11214
rect 14810 11121 14844 11137
rect 14810 8729 14844 8745
rect 14632 8652 14648 8686
rect 14748 8652 14764 8686
rect 14890 8652 14906 8686
rect 15006 8652 15022 8686
rect 15060 8532 15110 11333
rect 15576 8532 15626 11333
rect 16092 8532 16142 11333
rect 16180 11180 16196 11214
rect 16296 11180 16312 11214
rect 16438 11180 16454 11214
rect 16554 11180 16570 11214
rect 16358 11121 16392 11137
rect 16358 8729 16392 8745
rect 16180 8652 16196 8686
rect 16296 8652 16312 8686
rect 16438 8652 16454 8686
rect 16554 8652 16570 8686
rect 16608 8532 16658 11333
rect 16696 11180 16712 11214
rect 16812 11180 16828 11214
rect 16954 11180 16970 11214
rect 17070 11180 17086 11214
rect 16874 11121 16908 11137
rect 16874 8729 16908 8745
rect 16696 8652 16712 8686
rect 16812 8652 16828 8686
rect 16954 8652 16970 8686
rect 17070 8652 17086 8686
rect 17124 8532 17174 11333
rect 17212 11180 17228 11214
rect 17328 11180 17344 11214
rect 17470 11180 17486 11214
rect 17586 11180 17602 11214
rect 17390 11121 17424 11137
rect 17390 8729 17424 8745
rect 17212 8652 17228 8686
rect 17328 8652 17344 8686
rect 17470 8652 17486 8686
rect 17586 8652 17602 8686
rect 17640 8532 17690 11333
rect 18156 8532 18206 11333
rect 18672 8532 18722 11333
rect 18760 11180 18776 11214
rect 18876 11180 18892 11214
rect 19018 11180 19034 11214
rect 19134 11180 19150 11214
rect 18938 11121 18972 11137
rect 18938 8729 18972 8745
rect 18760 8652 18776 8686
rect 18876 8652 18892 8686
rect 19018 8652 19034 8686
rect 19134 8652 19150 8686
rect 19188 8532 19238 11333
rect 19276 11180 19292 11214
rect 19392 11180 19408 11214
rect 19534 11180 19550 11214
rect 19650 11180 19666 11214
rect 19454 11121 19488 11137
rect 19454 8729 19488 8745
rect 19276 8652 19292 8686
rect 19392 8652 19408 8686
rect 19534 8652 19550 8686
rect 19650 8652 19666 8686
rect 19704 8532 19754 11333
rect 20220 8532 20270 11333
rect 20308 11180 20324 11214
rect 20424 11180 20440 11214
rect 20566 11180 20582 11214
rect 20682 11180 20698 11214
rect 20486 11121 20520 11137
rect 20486 8729 20520 8745
rect 20308 8652 20324 8686
rect 20424 8652 20440 8686
rect 20566 8652 20582 8686
rect 20682 8652 20698 8686
rect 20736 8532 20786 11333
rect 21252 8532 21302 11333
rect 21590 10841 33411 11333
rect 21590 10672 22797 10841
rect 22990 10702 23126 10841
rect 24798 10704 25190 10841
rect 28410 10704 28802 10841
rect 30474 10704 30866 10841
rect 21590 9858 22954 10672
rect 21590 9666 22797 9858
rect 24968 9824 25018 10704
rect 28580 9824 28630 10704
rect 30644 9824 30694 10704
rect 32536 10700 32674 10841
rect 32844 10670 33411 10841
rect 32710 9856 33411 10670
rect 22990 9666 23126 9824
rect 24798 9666 25190 9824
rect 28410 9666 28802 9824
rect 30474 9666 30866 9824
rect 32538 9666 32672 9824
rect 32844 9678 33411 9856
rect 32812 9666 33411 9678
rect 21590 8876 33411 9666
rect 21590 8532 24212 8876
rect 9052 8055 24212 8532
rect 9052 8052 11358 8055
rect 11416 8052 24212 8055
rect 9052 8045 24212 8052
rect 4400 7456 4818 7624
rect 9052 7456 11686 8045
rect 16452 7864 16848 8045
rect 1162 6810 11686 7456
rect 1162 5310 3226 6810
rect 9379 6799 11686 6810
rect 9532 5310 11686 6799
rect 16616 5420 16682 7864
rect 1162 5096 2880 5310
rect 9867 5254 11686 5310
rect 16450 5258 16848 5420
rect 13256 5254 18299 5258
rect 9867 5250 18299 5254
rect 21612 5250 24212 8045
rect 9867 5102 24212 5250
rect 1162 3609 3220 5096
rect 9532 4690 24212 5102
rect 9532 3609 13844 4690
rect 15510 4522 15910 4690
rect 16802 4682 24212 4690
rect 15686 3616 15736 4522
rect 1162 3448 13844 3609
rect 15512 3448 15916 3616
rect 16802 3490 18640 4682
rect 19782 3490 20266 4682
rect 20730 3490 20784 4682
rect 21248 3502 24212 4682
rect 21248 3501 24285 3502
rect 24676 3501 24726 8876
rect 25192 3501 25242 8876
rect 25708 3501 25758 8876
rect 26224 3501 26274 8876
rect 26740 3501 26790 8876
rect 27256 3501 27306 8876
rect 27772 3501 27822 8876
rect 28288 3501 28338 8876
rect 28804 3501 28854 8876
rect 29320 3501 29370 8876
rect 29836 3501 29886 8876
rect 30352 3501 30402 8876
rect 30868 3501 30918 8876
rect 31384 3501 31434 8876
rect 31900 3501 31950 8876
rect 32420 3501 33411 8876
rect 21248 3490 33411 3501
rect 16802 3448 33411 3490
rect 1162 3442 33411 3448
rect -1704 3348 33411 3442
rect -3164 3342 33411 3348
rect -3742 3148 33411 3342
rect 33445 3466 33447 9678
rect -3776 3122 33445 3148
rect -3776 3088 -3716 3122
rect 33385 3088 33445 3122
rect -6420 2667 -3666 2796
rect -6426 2651 -3666 2667
rect -6346 2642 -3666 2651
rect -6346 2638 -4858 2642
rect -6346 2636 -6048 2638
rect -6346 -3658 -6058 2636
rect -5754 -3652 -4858 2638
rect -4564 2598 -3666 2642
rect -4564 2596 -2510 2598
rect -4564 2560 -2828 2596
rect -2776 2560 -2510 2596
rect -2460 2560 33460 2598
rect -4564 2558 -3004 2560
rect -4564 1806 -3662 2558
rect -3270 2452 -3004 2558
rect -3270 2418 -3060 2452
rect -3024 2420 -3004 2452
rect -2276 2556 33460 2560
rect -2276 2452 -2024 2556
rect -3024 2418 -3014 2420
rect -3270 2380 -3014 2418
rect -3406 2368 -3014 2380
rect -3406 1992 -3136 2368
rect -3102 1992 -3014 2368
rect -3406 1980 -3014 1992
rect -3270 1942 -3014 1980
rect -3270 1908 -3060 1942
rect -3024 1940 -3014 1942
rect -2276 2418 -2270 2452
rect -2230 2418 -2024 2452
rect -2276 2378 -2024 2418
rect -1628 2502 33460 2556
rect -1628 2414 33295 2502
rect -2276 2368 -1882 2378
rect -2276 1992 -2188 2368
rect -2154 1992 -1882 2368
rect -2276 1982 -1882 1992
rect -1628 2234 6476 2414
rect 6658 2252 6800 2414
rect 13108 2252 13248 2414
rect 13440 2240 33295 2414
rect -2276 1942 -2024 1982
rect -3024 1908 -3004 1940
rect -3270 1806 -3004 1908
rect -2276 1908 -2270 1942
rect -2230 1908 -2024 1942
rect -2276 1806 -2024 1908
rect -4564 1800 -2024 1806
rect -1628 1800 6624 2234
rect 13440 2230 14060 2240
rect -4564 1618 6624 1800
rect 13280 2064 14060 2230
rect 14258 2088 14400 2240
rect 16064 2088 16462 2240
rect 17356 2090 17494 2240
rect 13280 1654 14232 2064
rect -4564 1534 6480 1618
rect 13280 1614 14060 1654
rect 16240 1634 16288 2088
rect 17680 2066 18160 2240
rect 18358 2090 18496 2240
rect 19646 2080 20130 2240
rect 17680 2064 18324 2066
rect 17530 1654 18324 2064
rect 17680 1652 18324 1654
rect -4564 1364 -3018 1534
rect -2838 1390 -2706 1534
rect -4564 -248 -2876 1364
rect -4564 -420 -3018 -248
rect -2840 -420 -2704 -274
rect -2410 -420 -2360 1534
rect -1894 -420 -1844 1534
rect -1378 -420 -1328 1534
rect -862 -420 -812 1534
rect -346 -420 -296 1534
rect 170 -420 220 1534
rect 686 -420 736 1534
rect 1202 -420 1252 1534
rect 1548 1390 1680 1534
rect 1860 1458 6480 1534
rect 6654 1458 6798 1592
rect 1860 1402 6802 1458
rect 13108 1448 13248 1592
rect 13440 1480 14060 1614
rect 14262 1480 14398 1630
rect 16062 1480 16468 1634
rect 17358 1480 17496 1630
rect 17680 1480 18160 1652
rect 19822 1636 19872 2080
rect 20080 1636 20130 2080
rect 18360 1480 18498 1628
rect 19650 1480 20130 1636
rect 20596 1480 20646 2240
rect 21112 2090 21334 2240
rect 21112 1624 21162 2090
rect 21520 2064 33295 2240
rect 21370 1984 33295 2064
rect 21370 1814 22554 1984
rect 22734 1838 22866 1984
rect 21370 1650 22694 1814
rect 21112 1480 21336 1624
rect 21520 1480 22694 1650
rect 13440 1448 22694 1480
rect 13108 1412 22694 1448
rect 1860 1362 6480 1402
rect 1718 1246 6480 1362
rect 6654 1268 6798 1402
rect 13110 1268 13248 1412
rect 13440 1246 22694 1412
rect 1718 840 6628 1246
rect 1718 664 2560 840
rect 2740 694 2816 840
rect 4164 696 4236 840
rect 1718 -246 2722 664
rect 4420 658 6628 840
rect 4256 630 6628 658
rect 9924 630 9980 1246
rect 13282 660 22694 1246
rect 13282 630 14080 660
rect 4256 440 6480 630
rect 6658 440 6796 612
rect 13110 440 13248 608
rect 13440 462 14080 630
rect 14262 490 14394 660
rect 17616 488 18006 660
rect 21228 490 21360 660
rect 13440 440 14222 462
rect 4256 40 14222 440
rect 4256 -138 5460 40
rect 5662 -112 5794 40
rect 6952 -110 7342 40
rect 4256 -242 5622 -138
rect 1860 -248 2722 -246
rect 1548 -420 1680 -272
rect 1860 -420 2560 -248
rect 2740 -420 2816 -278
rect 4164 -420 4236 -280
rect 4420 -420 5622 -242
rect -4564 -512 5622 -420
rect -4564 -1296 -3896 -512
rect -3472 -1046 5622 -512
rect -3472 -1060 5480 -1046
rect -3472 -1228 -3020 -1060
rect -2800 -1210 -2544 -1060
rect -1426 -1208 -1170 -1060
rect -3472 -1296 -2880 -1228
rect -4564 -1654 -2880 -1296
rect -4564 -1820 -3020 -1654
rect -2804 -1820 -2542 -1676
rect -1428 -1820 -1172 -1666
rect -1092 -1820 -1046 -1060
rect -968 -1210 -712 -1060
rect 4072 -1212 4326 -1060
rect 4540 -1220 5480 -1060
rect 5662 -1220 5794 -1072
rect 6952 -1074 7084 -1072
rect 7124 -1074 7170 -110
rect 8496 -112 8898 40
rect 13142 -110 13278 40
rect 8670 -1072 8722 -112
rect 13440 -136 14222 40
rect 13314 -746 14222 -136
rect 17788 -746 17834 488
rect 21560 462 22694 660
rect 21400 -196 22694 462
rect 21400 -368 22554 -196
rect 22734 -368 22866 -220
rect 22906 -368 22952 1984
rect 23422 -368 23468 1984
rect 23938 -368 23984 1984
rect 24454 -368 24500 1984
rect 24970 -368 25016 1984
rect 25486 -368 25532 1984
rect 26002 -368 26048 1984
rect 26518 -368 26564 1984
rect 27034 -368 27080 1984
rect 27550 -368 27596 1984
rect 28066 -368 28112 1984
rect 28582 -368 28628 1984
rect 29098 -368 29144 1984
rect 29614 -368 29660 1984
rect 30130 -368 30176 1984
rect 30646 -368 30692 1984
rect 31162 -368 31208 1984
rect 31246 1838 31382 1984
rect 31560 1814 33295 1984
rect 31420 1670 33295 1814
rect 31420 -196 31920 1670
rect 31248 -368 31380 -220
rect 31560 -368 31920 -196
rect 21400 -386 31920 -368
rect 21400 -396 31982 -386
rect 33010 -396 33295 1670
rect 21400 -746 33295 -396
rect 13314 -920 14080 -746
rect 14262 -920 14394 -772
rect 17616 -920 18006 -746
rect 21228 -920 21360 -774
rect 21560 -920 33295 -746
rect 13314 -940 33295 -920
rect 13314 -1054 22160 -940
rect 6952 -1220 7342 -1074
rect 8500 -1220 8890 -1072
rect 13142 -1220 13282 -1070
rect 13440 -1136 22160 -1054
rect 22360 -1110 22496 -940
rect 23134 -1112 23528 -940
rect 25972 -942 26108 -940
rect 26144 -942 26194 -940
rect 26230 -1112 26624 -940
rect 13440 -1220 22324 -1136
rect 4540 -1236 22324 -1220
rect 4408 -1460 22324 -1236
rect 4408 -1638 14080 -1460
rect 14262 -1612 14394 -1460
rect 4408 -1646 14222 -1638
rect -968 -1820 -712 -1666
rect 4072 -1820 4326 -1672
rect 4540 -1760 14222 -1646
rect 4540 -1820 6480 -1760
rect -4564 -1938 6480 -1820
rect 6662 -1910 6794 -1760
rect -4564 -2196 6624 -1938
rect -4564 -2976 -3902 -2196
rect -3474 -2260 6624 -2196
rect -3474 -2436 -3020 -2260
rect -2792 -2400 -2546 -2260
rect -3474 -2842 -2888 -2436
rect -3474 -2976 -3020 -2842
rect -4564 -3020 -3020 -2976
rect -2800 -3020 -2548 -2886
rect -2008 -3020 -1962 -2260
rect -1092 -3020 -1046 -2260
rect -176 -3020 -130 -2260
rect 266 -3020 286 -3018
rect 740 -3020 786 -2260
rect 1656 -3020 1702 -2260
rect 2572 -3020 2618 -2260
rect 3160 -2400 3412 -2260
rect 3620 -2360 6624 -2260
rect 3620 -2442 4180 -2360
rect 3494 -2538 4180 -2442
rect 3494 -2840 4324 -2538
rect 3620 -2846 4324 -2840
rect 4680 -2846 6624 -2360
rect 3154 -3020 3406 -2882
rect 3620 -3020 4180 -2846
rect 4680 -3020 6480 -2846
rect -4564 -3040 6480 -3020
rect 6662 -3040 6794 -2872
rect 7090 -3040 7140 -1760
rect 7606 -3040 7656 -1760
rect 8122 -3040 8172 -1760
rect 8638 -3040 8688 -1760
rect 9154 -3040 9204 -1760
rect 9670 -3040 9720 -1760
rect 10186 -3040 10236 -1760
rect 10702 -3040 10752 -1760
rect 11218 -3040 11268 -1760
rect 11734 -3040 11784 -1760
rect 12250 -3040 12300 -1760
rect 12766 -3040 12816 -1760
rect 13112 -1910 13244 -1760
rect 13440 -1938 14222 -1760
rect 13284 -2846 14222 -1938
rect 13112 -3040 13244 -2872
rect 13440 -3040 14080 -2846
rect 14262 -3040 14394 -2872
rect 14432 -3040 14482 -1460
rect 14948 -3040 14998 -1460
rect 15464 -3040 15514 -1460
rect 15980 -3040 16030 -1460
rect 16496 -3040 16546 -1460
rect 17012 -3040 17062 -1460
rect 17528 -3040 17578 -1460
rect 18044 -3040 18094 -1460
rect 18560 -3040 18610 -1460
rect 19076 -3040 19126 -1460
rect 19592 -3040 19642 -1460
rect 20108 -3040 20158 -1460
rect 20624 -3040 20674 -1460
rect 20712 -1610 20844 -1460
rect 21040 -1548 22324 -1460
rect 21040 -1638 22160 -1548
rect 23306 -1572 23356 -1112
rect 26402 -1572 26452 -1112
rect 29324 -1114 29720 -940
rect 32422 -1114 32558 -940
rect 29498 -1570 29548 -1114
rect 32740 -1134 33295 -940
rect 32596 -1548 33295 -1134
rect 20882 -1720 22160 -1638
rect 22362 -1720 22494 -1574
rect 23134 -1720 23528 -1572
rect 20882 -1740 23660 -1720
rect 26230 -1740 26628 -1572
rect 29326 -1740 29720 -1570
rect 32422 -1740 32560 -1570
rect 32740 -1740 33295 -1548
rect 20882 -2180 33295 -1740
rect 20882 -2374 22180 -2180
rect 22374 -2330 22500 -2180
rect 20882 -2772 22328 -2374
rect 20882 -2846 22180 -2772
rect 20712 -3040 20844 -2870
rect 21040 -2962 22180 -2846
rect 22378 -2962 22504 -2806
rect 22800 -2962 22850 -2180
rect 23316 -2962 23366 -2180
rect 23832 -2962 23882 -2180
rect 24176 -2342 24568 -2180
rect 24352 -2806 24394 -2342
rect 24178 -2962 24570 -2806
rect 24866 -2962 24912 -2180
rect 25382 -2962 25428 -2180
rect 25898 -2962 25944 -2180
rect 26416 -2962 26462 -2180
rect 26932 -2962 26974 -2180
rect 27446 -2962 27488 -2180
rect 27960 -2962 28008 -2180
rect 28476 -2962 28526 -2180
rect 28992 -2962 29042 -2180
rect 29508 -2962 29558 -2180
rect 29854 -2342 30246 -2180
rect 30028 -2800 30070 -2342
rect 29854 -2962 30244 -2800
rect 30540 -2962 30590 -2180
rect 31056 -2962 31106 -2180
rect 31572 -2962 31622 -2180
rect 31918 -2316 32048 -2180
rect 32244 -2372 33295 -2180
rect 32090 -2776 33295 -2372
rect 31918 -2962 32048 -2814
rect 32244 -2962 33295 -2776
rect 21040 -3040 33295 -2962
rect -4564 -3652 33295 -3040
rect -5754 -3656 33295 -3652
rect -5764 -3658 33295 -3656
rect -6346 -4728 33295 -3658
rect -6346 -5124 -4414 -4728
rect -6426 -5140 -4414 -5124
rect -6410 -5410 -4414 -5140
rect 33248 -4863 33295 -4728
rect 33427 -3637 33460 2502
rect 33248 -4879 33427 -4863
rect -6410 -5589 -6206 -5410
rect -6410 -5596 -4414 -5589
rect 33248 -5596 33426 -4879
rect -6410 -5622 33426 -5596
rect -7724 -6803 -7594 -6456
rect -7229 -6476 -7195 -6450
rect 50952 -6476 50986 -6450
rect -7229 -6510 -7169 -6476
rect 50926 -6510 50986 -6476
rect 51264 15918 51330 16138
rect 51327 15916 51330 15918
rect 51264 -6680 51327 -6670
rect 51264 -6686 51332 -6680
rect 51268 -6798 51332 -6686
rect 51038 -6803 51340 -6798
rect -7724 -6916 -7686 -6803
rect -7702 -6929 -7686 -6916
rect 51106 -6926 51340 -6803
rect 51106 -6929 51122 -6926
<< viali >>
rect -9948 4985 -9418 5157
rect -9960 3449 -9336 3623
rect -3384 14434 33104 15092
rect -2992 4702 -2936 4744
rect -2680 4700 -2624 4742
rect -2362 4706 -2306 4748
rect -2828 2560 -2776 2596
rect -2510 2560 -2460 2598
rect -3136 1992 -3102 2368
rect -2270 2418 -2230 2452
rect -2188 1992 -2154 2368
rect -2270 1908 -2230 1942
rect -4414 -5410 33248 -4728
rect -4414 -5589 33230 -5410
rect 33230 -5589 33248 -5410
rect -4414 -5596 33248 -5589
<< metal1 >>
rect -6482 15092 33382 15434
rect -6482 14434 -3384 15092
rect 33104 14434 33382 15092
rect -6482 14312 33382 14434
rect -4182 14100 -4121 14106
rect -5414 13786 -5330 13802
rect -5414 13702 -5332 13786
rect -5248 13702 -5242 13786
rect -9960 5157 -9406 5163
rect -9960 4985 -9948 5157
rect -9418 4985 -9406 5157
rect -9960 4979 -9406 4985
rect -5614 5086 -5550 5092
rect -9426 4859 -9256 4893
rect -9970 4219 -9652 4389
rect -9426 4366 -9392 4859
rect -8615 4857 -8442 4895
rect -9258 4557 -9031 4619
rect -9426 4332 -9259 4366
rect -9305 4219 -9271 4332
rect -9093 4266 -9031 4557
rect -8615 4368 -8577 4857
rect -8436 4531 -8230 4595
rect -8615 4330 -8453 4368
rect -8491 4266 -8453 4330
rect -9970 4173 -9270 4219
rect -9093 4204 -8453 4266
rect -9970 4059 -9652 4173
rect -9305 4056 -9271 4173
rect -9435 4022 -9271 4056
rect -9435 3740 -9401 4022
rect -9093 3916 -9031 4204
rect -9267 3854 -9031 3916
rect -9435 3706 -9267 3740
rect -9972 3623 -9324 3629
rect -9972 3449 -9960 3623
rect -9336 3449 -9324 3623
rect -9972 3443 -9324 3449
rect -8903 3346 -8841 4204
rect -8491 4056 -8453 4204
rect -8639 4018 -8453 4056
rect -8294 4249 -8230 4531
rect -8294 4185 -8186 4249
rect -8122 4185 -8116 4249
rect -8639 3742 -8601 4018
rect -8294 3911 -8230 4185
rect -8442 3847 -8230 3911
rect -8639 3704 -8453 3742
rect -8903 3278 -8841 3284
rect -6000 2762 -5948 2768
rect -6000 2704 -5948 2710
rect -5996 -3524 -5952 2704
rect -5614 2258 -5550 5022
rect -5414 2762 -5330 13702
rect -4182 7694 -4121 14039
rect 23339 14100 23400 14106
rect -3947 13899 -3889 13905
rect -3947 7909 -3889 13841
rect -3771 13755 -3705 13761
rect -3771 8131 -3705 13689
rect -3561 13535 -3499 13541
rect -3561 8379 -3499 13473
rect 17467 13535 17529 13541
rect -3445 13399 -3387 13405
rect -3445 8493 -3387 13341
rect 17191 13399 17249 13405
rect -3334 13266 -3266 13272
rect -3334 8606 -3266 13198
rect 16971 13265 17037 13271
rect -3208 13134 -3148 13140
rect -3208 8706 -3148 13074
rect 11808 13014 11880 13020
rect 2782 12980 2834 12986
rect 2782 12922 2834 12928
rect 11554 12980 11606 12986
rect 11554 12922 11606 12928
rect -2916 12832 -2856 12838
rect -2916 12766 -2856 12772
rect 2186 12832 2246 12838
rect -3080 12632 -3008 12638
rect -3080 8974 -3008 12560
rect -3080 8896 -3008 8902
rect -2913 8809 -2859 12766
rect -610 12624 -560 12748
rect -780 12622 -392 12624
rect -94 12622 -44 12752
rect 2186 12642 2246 12772
rect -2334 12570 -2324 12622
rect -2200 12570 -2190 12622
rect -2076 12570 -2066 12622
rect -1942 12570 -1932 12622
rect -1818 12570 -1808 12622
rect -1684 12570 -1674 12622
rect -1560 12570 -1550 12622
rect -1426 12570 -1416 12622
rect -1302 12570 -1292 12622
rect -1168 12570 -1158 12622
rect -1044 12570 -1034 12622
rect -910 12570 -900 12622
rect -786 12570 -776 12622
rect -652 12570 -518 12622
rect -394 12570 -384 12622
rect -270 12570 -260 12622
rect -136 12570 -2 12622
rect 122 12570 132 12622
rect 246 12570 256 12622
rect 380 12570 390 12622
rect 504 12570 514 12622
rect 638 12570 648 12622
rect 762 12570 772 12622
rect 896 12570 906 12622
rect 1020 12570 1030 12622
rect 1154 12570 1164 12622
rect 1278 12570 1288 12622
rect 1412 12570 1422 12622
rect 1536 12570 1546 12622
rect 1670 12570 1680 12622
rect 2186 12576 2246 12582
rect -2324 9242 -2200 12570
rect -2158 9161 -2108 12538
rect -2066 9242 -1942 12570
rect -1808 9242 -1684 12570
rect -1642 9161 -1592 12538
rect -1550 9242 -1426 12570
rect -1292 9242 -1168 12570
rect -1126 9161 -1076 12538
rect -1034 9242 -910 12570
rect -780 12568 -392 12570
rect -776 9242 -652 12568
rect -610 9320 -560 12568
rect -518 9242 -394 12568
rect -260 9242 -136 12570
rect -94 9324 -44 12570
rect -2 9242 122 12570
rect 256 9242 380 12570
rect 424 9161 474 12538
rect 514 9242 638 12570
rect 772 9242 896 12570
rect 938 9161 988 12538
rect 1030 9242 1154 12570
rect 1288 9242 1412 12570
rect 1454 9183 1504 12538
rect 1546 9242 1670 12570
rect 2596 12516 2676 12522
rect 2418 9934 2470 9938
rect 2416 9932 2472 9934
rect 2416 9880 2418 9932
rect 2470 9880 2472 9932
rect 2256 9802 2308 9808
rect 2256 9744 2308 9750
rect 1441 9161 1535 9183
rect -2158 9111 1535 9161
rect -2158 9110 -2108 9111
rect -1642 9110 -1592 9111
rect -1126 9110 -1076 9111
rect 424 9110 474 9111
rect 938 9110 988 9111
rect -2913 8749 -2859 8755
rect -986 8976 -930 8982
rect -3208 8640 -3148 8646
rect -3334 8532 -3266 8538
rect -3445 8429 -3387 8435
rect -3561 8311 -3499 8317
rect -1607 8131 -1541 8137
rect -3777 8065 -3771 8131
rect -3705 8065 -3699 8131
rect -3947 7845 -3889 7851
rect -1755 7909 -1697 7915
rect -4182 7627 -4121 7633
rect -1918 7694 -1857 7700
rect -3812 6308 -3748 6314
rect -3812 5086 -3748 6244
rect -1918 6095 -1857 7633
rect -1755 6895 -1697 7851
rect -1607 7075 -1541 8065
rect -1607 7003 -1541 7009
rect -1755 6831 -1697 6837
rect -1581 6895 -1523 6901
rect -1924 6034 -1918 6095
rect -1857 6034 -1851 6095
rect -1760 6094 -1700 6100
rect -3172 5960 -3162 5964
rect -3812 5016 -3748 5022
rect -3667 5902 -3162 5960
rect -3667 4437 -3609 5902
rect -3172 5900 -3162 5902
rect -3076 5960 -3066 5964
rect -3076 5902 -3064 5960
rect -3076 5900 -3066 5902
rect -3392 5784 -3328 5830
rect -3234 5784 -3170 5830
rect -3462 4943 -3416 5743
rect -3374 4902 -3342 5784
rect -3304 4943 -3258 5743
rect -3222 4904 -3192 5784
rect -3140 5743 -3106 5900
rect -2208 5892 -2198 5958
rect -2140 5892 -2130 5958
rect -3076 5784 -3012 5830
rect -3146 4943 -3100 5743
rect -3058 4904 -3026 5784
rect -2932 5778 -2922 5836
rect -2374 5778 -2364 5836
rect -2286 5784 -2222 5830
rect -2982 5743 -2948 5748
rect -2988 4943 -2942 5743
rect -3392 4856 -3328 4902
rect -3264 4838 -3254 4904
rect -3022 4838 -3012 4904
rect -2982 4750 -2948 4943
rect -2902 4902 -2870 5778
rect -2830 4934 -2784 5748
rect -2918 4856 -2854 4902
rect -3004 4744 -2924 4750
rect -3004 4702 -2992 4744
rect -2936 4702 -2924 4744
rect -2826 4728 -2788 4934
rect -2744 4902 -2712 5778
rect -2666 5743 -2632 5748
rect -2672 4943 -2626 5743
rect -2760 4856 -2696 4902
rect -2666 4748 -2632 4943
rect -2584 4902 -2552 5778
rect -2514 4943 -2468 5743
rect -2602 4856 -2538 4902
rect -2508 4764 -2474 4943
rect -2430 4902 -2398 5778
rect -2350 5743 -2316 5748
rect -2356 4943 -2310 5743
rect -2444 4856 -2380 4902
rect -2692 4742 -2612 4748
rect -3004 4696 -2924 4702
rect -2854 4664 -2844 4728
rect -2768 4664 -2758 4728
rect -2692 4700 -2680 4742
rect -2624 4700 -2612 4742
rect -2512 4728 -2464 4764
rect -2350 4754 -2316 4943
rect -2270 4912 -2238 5784
rect -2192 5743 -2158 5892
rect -2128 5784 -2064 5830
rect -1970 5784 -1906 5830
rect -2198 4943 -2152 5743
rect -2110 4912 -2078 5784
rect -2040 4943 -1994 5743
rect -2284 4902 -2274 4912
rect -2286 4856 -2274 4902
rect -2284 4846 -2274 4856
rect -2042 4846 -2032 4912
rect -1954 4902 -1922 5784
rect -1882 4943 -1836 5743
rect -1970 4856 -1906 4902
rect -2374 4748 -2294 4754
rect -2692 4694 -2612 4700
rect -2538 4664 -2528 4728
rect -2452 4664 -2442 4728
rect -2374 4706 -2362 4748
rect -2306 4706 -2294 4748
rect -2374 4700 -2294 4706
rect -3667 4379 -3337 4437
rect -2512 4432 -2464 4664
rect -1760 4660 -1700 6034
rect -1581 5867 -1523 6837
rect -1581 5803 -1523 5809
rect -1760 4594 -1700 4600
rect -2512 4384 -1890 4432
rect -4028 4252 -3964 4258
rect -4210 3354 -4138 3360
rect -4562 3068 -4490 3074
rect -5178 2876 -5126 2882
rect -5178 2818 -5126 2824
rect -5414 2710 -5398 2762
rect -5346 2710 -5330 2762
rect -5414 2694 -5330 2710
rect -5904 2194 -5550 2258
rect -5910 1460 -5864 1654
rect -5173 1463 -5131 2818
rect -4798 2762 -4746 2768
rect -4798 2704 -4746 2710
rect -5910 1457 -5790 1460
rect -5178 1457 -5126 1463
rect -5910 1405 -5846 1457
rect -5794 1405 -5788 1457
rect -5910 1404 -5790 1405
rect -5910 1250 -5864 1404
rect -5178 1399 -5126 1405
rect -5912 670 -5864 868
rect -5137 670 -5079 676
rect -5912 612 -5889 670
rect -5831 612 -5780 670
rect -5912 464 -5864 612
rect -5906 -126 -5858 84
rect -5906 -128 -5792 -126
rect -5906 -180 -5850 -128
rect -5798 -180 -5792 -128
rect -5236 -128 -5184 -122
rect -5906 -318 -5858 -180
rect -5236 -186 -5184 -180
rect -5902 -874 -5814 -706
rect -5386 -874 -5279 -868
rect -5902 -960 -5803 -874
rect -5717 -960 -5658 -874
rect -5386 -960 -5365 -874
rect -5902 -1100 -5814 -960
rect -5386 -966 -5279 -960
rect -5902 -1700 -5864 -1490
rect -5902 -1709 -5822 -1700
rect -5902 -1761 -5880 -1709
rect -5828 -1761 -5822 -1709
rect -5902 -1768 -5822 -1761
rect -5486 -1704 -5410 -1696
rect -5486 -1766 -5479 -1704
rect -5417 -1766 -5410 -1704
rect -5902 -1890 -5864 -1768
rect -5486 -1774 -5410 -1766
rect -5904 -2470 -5860 -2268
rect -5904 -2481 -5814 -2470
rect -5904 -2533 -5875 -2481
rect -5823 -2533 -5814 -2481
rect -5904 -2544 -5814 -2533
rect -5584 -2481 -5532 -2475
rect -5584 -2539 -5532 -2533
rect -5904 -2678 -5860 -2544
rect -5900 -3285 -5868 -3050
rect -5690 -3285 -5638 -3279
rect -5900 -3337 -5876 -3285
rect -5824 -3337 -5818 -3285
rect -5900 -3470 -5868 -3337
rect -5690 -3343 -5638 -3337
rect -5994 -3534 -5962 -3524
rect -5687 -3920 -5641 -3343
rect -5579 -3818 -5537 -2539
rect -5471 -3704 -5425 -1774
rect -5474 -3710 -5422 -3704
rect -5474 -3768 -5422 -3762
rect -5584 -3824 -5532 -3818
rect -5584 -3882 -5532 -3876
rect -5696 -3972 -5690 -3920
rect -5638 -3972 -5632 -3920
rect -5346 -4020 -5294 -966
rect -5358 -4029 -5285 -4020
rect -5358 -4108 -5285 -4102
rect -5229 -4210 -5191 -186
rect -5236 -4216 -5184 -4210
rect -5236 -4274 -5184 -4268
rect -5137 -4341 -5079 612
rect -4791 -3529 -4752 2704
rect -4562 2296 -4490 2996
rect -4430 2876 -4378 2882
rect -4430 2818 -4378 2824
rect -4702 2224 -4490 2296
rect -4700 1446 -4658 1660
rect -4425 1596 -4383 2818
rect -4210 1952 -4138 3282
rect -4028 2480 -3964 4188
rect -3484 4016 -3420 4210
rect -3634 3972 -3420 4016
rect -3864 2850 -3812 2856
rect -3864 2792 -3812 2798
rect -4028 2410 -3964 2416
rect -4210 1874 -4138 1880
rect -4430 1590 -4378 1596
rect -4430 1532 -4378 1538
rect -3862 1454 -3814 2792
rect -3634 2762 -3590 3972
rect -3484 3540 -3420 3972
rect -3383 3351 -3349 4379
rect -3676 2710 -3670 2762
rect -3618 2710 -3590 2762
rect -3634 2380 -3590 2710
rect -3484 3317 -3349 3351
rect -1929 3367 -1895 4384
rect -1846 3922 -1642 3978
rect -1929 3333 -1808 3367
rect -3484 2672 -3450 3317
rect -3502 2666 -3450 2672
rect -3502 2608 -3450 2614
rect -2671 2666 -2619 2672
rect -2671 2608 -2619 2614
rect -3634 2306 -3524 2380
rect -3598 1980 -3524 2306
rect -3484 1910 -3450 2608
rect -2840 2596 -2764 2602
rect -2840 2560 -2828 2596
rect -2776 2560 -2764 2596
rect -2840 2550 -2764 2560
rect -3072 2452 -3008 2458
rect -3072 2418 -3060 2452
rect -3024 2418 -3008 2452
rect -2924 2418 -2914 2470
rect -2862 2458 -2852 2470
rect -2862 2418 -2850 2458
rect -3072 2412 -3008 2418
rect -2914 2412 -2850 2418
rect -3142 2368 -3096 2380
rect -3142 1992 -3136 2368
rect -3102 1992 -3096 2368
rect -3142 1980 -3096 1992
rect -3052 1948 -3024 2412
rect -2978 2380 -2944 2382
rect -2984 1980 -2938 2380
rect -3072 1942 -3008 1948
rect -3072 1908 -3060 1942
rect -3024 1908 -3008 1942
rect -3072 1902 -3008 1908
rect -2978 1830 -2944 1980
rect -2898 1948 -2870 2412
rect -2820 2380 -2786 2550
rect -2756 2412 -2692 2458
rect -2826 1980 -2780 2380
rect -2738 1948 -2710 2412
rect -2662 2380 -2628 2608
rect -2522 2598 -2448 2604
rect -2522 2560 -2510 2598
rect -2460 2560 -2448 2598
rect -2522 2548 -2448 2560
rect -2598 2412 -2534 2458
rect -2668 1980 -2622 2380
rect -2662 1976 -2628 1980
rect -2580 1948 -2552 2412
rect -2504 2380 -2470 2548
rect -2438 2458 -2428 2470
rect -2440 2418 -2428 2458
rect -2376 2418 -2366 2470
rect -2282 2452 -2218 2458
rect -2282 2418 -2270 2452
rect -2230 2418 -2218 2452
rect -2440 2412 -2376 2418
rect -2282 2412 -2218 2418
rect -2510 1980 -2464 2380
rect -2424 1948 -2396 2412
rect -2346 2380 -2312 2382
rect -2352 1980 -2306 2380
rect -2914 1902 -2850 1948
rect -2756 1942 -2692 1948
rect -2766 1890 -2756 1942
rect -2704 1902 -2692 1942
rect -2598 1942 -2534 1948
rect -2598 1902 -2586 1942
rect -2704 1890 -2694 1902
rect -2596 1890 -2586 1902
rect -2534 1890 -2524 1942
rect -2440 1902 -2376 1948
rect -2346 1830 -2312 1980
rect -2266 1948 -2230 2412
rect -2194 2368 -2148 2380
rect -2194 1992 -2188 2368
rect -2154 1992 -2148 2368
rect -2194 1980 -2148 1992
rect -1842 1981 -1808 3333
rect -1698 3324 -1642 3922
rect -1229 3330 -1183 8137
rect -1140 7664 -1042 8046
rect -986 7664 -930 8920
rect 322 8706 382 8712
rect -533 8493 -475 8499
rect -1140 7608 -930 7664
rect -653 8379 -591 8385
rect -1140 7250 -1042 7608
rect -913 7075 -847 7081
rect -1146 6476 -1034 6844
rect -913 6476 -847 7009
rect -1146 6410 -847 6476
rect -1146 6034 -1034 6410
rect -653 6306 -591 8317
rect -533 7738 -475 8435
rect -410 7738 -358 8054
rect -533 7680 -358 7738
rect -410 7238 -358 7680
rect -420 6306 -360 6846
rect -660 6230 -360 6306
rect -420 6030 -360 6230
rect -601 5809 -595 5867
rect -537 5809 -531 5867
rect -1142 4942 -1072 5642
rect -595 5308 -537 5809
rect -422 5308 -356 5642
rect -595 5250 -356 5308
rect -1142 4882 -986 4942
rect -926 4882 -920 4942
rect -1142 4828 -1072 4882
rect -422 4826 -356 5250
rect -1154 3756 -1052 4446
rect -472 3768 -356 4438
rect -1154 3698 -937 3756
rect -1154 3624 -1052 3698
rect -1234 3324 -1178 3330
rect -1698 3268 -1636 3324
rect -1580 3268 -1574 3324
rect -1698 2958 -1642 3268
rect -1234 3262 -1178 3268
rect -1708 2904 -1698 2958
rect -1644 2904 -1634 2958
rect -1698 2382 -1642 2904
rect -1500 2850 -1448 2856
rect -1500 2792 -1448 2798
rect -1768 2278 -1642 2382
rect -2282 1942 -2218 1948
rect -2282 1908 -2270 1942
rect -2230 1908 -2218 1942
rect -2282 1902 -2218 1908
rect -1845 1830 -1807 1981
rect -1768 1978 -1684 2278
rect -1498 1952 -1450 2792
rect -995 2703 -937 3698
rect -590 3720 -356 3768
rect -590 3168 -542 3720
rect -472 3622 -356 3720
rect -325 3330 -287 8129
rect 101 3330 144 8133
rect 180 7704 242 8046
rect 322 7704 382 8646
rect 180 7644 382 7704
rect 433 8607 503 8613
rect 180 7242 242 7644
rect 178 6388 244 6840
rect 433 6388 503 8537
rect 791 8541 853 8547
rect 791 7650 853 8479
rect 936 7650 1024 8044
rect 791 7588 1024 7650
rect 936 7244 1024 7588
rect 796 7068 857 7074
rect 796 6428 857 7007
rect 968 6428 1028 6846
rect 178 6314 505 6388
rect 790 6356 1028 6428
rect 178 6044 244 6314
rect 968 6028 1028 6356
rect 793 5865 851 5871
rect 180 4932 260 5638
rect 793 5234 851 5807
rect 928 5234 1028 5632
rect 779 5148 1028 5234
rect 180 4866 561 4932
rect 180 4838 260 4866
rect 180 3716 240 4444
rect 180 3652 428 3716
rect 180 3630 240 3652
rect 364 3522 428 3652
rect 364 3452 428 3458
rect -334 3324 -278 3330
rect -334 3262 -278 3268
rect 94 3324 150 3330
rect 94 3262 150 3268
rect -592 3162 -540 3168
rect -592 3104 -540 3110
rect 495 2797 561 4866
rect 928 4834 1028 5148
rect 806 4668 862 4674
rect 806 4020 862 4612
rect 974 4020 1024 4434
rect 806 3964 1024 4020
rect 974 3626 1024 3964
rect 1062 3330 1106 8128
rect 1441 7387 1535 9111
rect 1894 8974 1966 8980
rect 1441 7287 1535 7293
rect 1689 8809 1743 8815
rect 1056 3324 1112 3330
rect 1056 3262 1112 3268
rect 1525 3277 1583 3283
rect 495 2725 561 2731
rect -995 2639 -937 2645
rect -1500 1946 -1448 1952
rect -1500 1888 -1448 1894
rect -2978 1792 -1807 1830
rect -3185 1717 -3127 1723
rect -3864 1448 -3812 1454
rect -4588 1446 -4582 1448
rect -4700 1398 -4582 1446
rect -4700 1254 -4658 1398
rect -4588 1396 -4582 1398
rect -4530 1396 -4524 1448
rect -3864 1390 -3812 1396
rect -4704 660 -4634 866
rect -3185 660 -3127 1659
rect 1525 1717 1583 3219
rect 1525 1653 1583 1659
rect -2913 1591 -2859 1596
rect -2576 1595 1418 1616
rect 1689 1595 1743 8755
rect 1894 1826 1966 8902
rect 1894 1748 1966 1754
rect 2090 8432 2166 8438
rect -2576 1591 1743 1595
rect -2913 1590 1743 1591
rect -2913 1538 -2524 1590
rect -2472 1574 1743 1590
rect -2472 1538 -2452 1574
rect -2913 1537 -2452 1538
rect -4704 602 -4621 660
rect -4563 602 -4557 660
rect -4704 472 -4634 602
rect -3185 596 -3127 602
rect -4694 -108 -4648 88
rect -4267 -108 -4213 -102
rect -4694 -162 -4672 -108
rect -4618 -162 -4612 -108
rect -4694 -312 -4648 -162
rect -4692 -792 -4640 -722
rect -4692 -844 -4634 -792
rect -4582 -844 -4576 -792
rect -4692 -1074 -4640 -844
rect -4685 -1625 -4623 -1505
rect -4685 -1863 -4623 -1687
rect -4416 -1958 -4351 -1952
rect -4416 -2445 -4351 -2023
rect -4700 -2510 -4351 -2445
rect -4698 -3184 -4664 -3062
rect -4698 -3190 -4581 -3184
rect -4698 -3300 -4691 -3190
rect -4698 -3306 -4581 -3300
rect -4698 -3450 -4664 -3306
rect -4788 -3532 -4756 -3529
rect -4267 -3543 -4213 -162
rect -3955 -447 -3881 -441
rect -4132 -792 -4080 -786
rect -4132 -3458 -4080 -844
rect -3955 -869 -3881 -521
rect -3241 -447 -3167 -441
rect -2668 -462 -2618 1364
rect -2576 -320 -2452 1537
rect -2318 -320 -2194 1574
rect -2152 -462 -2102 1364
rect -2060 -320 -1936 1574
rect -1802 -320 -1678 1574
rect -1636 -248 -1586 1574
rect -1544 -320 -1420 1574
rect -1286 -320 -1162 1574
rect -1120 -462 -1070 1364
rect -1028 -320 -904 1574
rect -770 -320 -646 1574
rect -604 -462 -554 1364
rect -512 -320 -388 1574
rect -254 -320 -130 1574
rect -88 -462 -38 1364
rect 4 -320 128 1574
rect 262 -320 386 1574
rect 428 -248 478 1574
rect 520 -320 644 1574
rect 778 -320 902 1574
rect 944 -462 994 1364
rect 1036 -320 1160 1574
rect 1294 1541 1743 1574
rect 1294 -320 1418 1541
rect 1460 -448 1510 1364
rect 1338 -462 1348 -448
rect -2668 -502 1348 -462
rect 1510 -502 1520 -448
rect -3750 -668 -3740 -588
rect -3636 -668 -3626 -588
rect -3790 -869 -3744 -700
rect -3955 -943 -3744 -869
rect -3790 -1100 -3744 -943
rect -3708 -1132 -3670 -668
rect -3632 -954 -3584 -700
rect -3241 -802 -3167 -521
rect -2346 -866 -2336 -812
rect -2092 -866 -2082 -812
rect -1888 -866 -1878 -812
rect -1634 -866 -1624 -812
rect -514 -866 -504 -812
rect -260 -866 -250 -812
rect -56 -866 -46 -812
rect 198 -866 208 -812
rect 402 -866 412 -812
rect 656 -866 666 -812
rect 860 -866 870 -812
rect 1114 -866 1124 -812
rect 1318 -866 1328 -812
rect 1572 -866 1582 -812
rect 1776 -866 1786 -812
rect 2030 -866 2040 -812
rect -3241 -882 -3167 -876
rect -3632 -960 -3436 -954
rect -3632 -1036 -3584 -960
rect -3458 -1036 -3436 -960
rect -3632 -1042 -3436 -1036
rect -3632 -1100 -3584 -1042
rect -3748 -1208 -3738 -1132
rect -3644 -1208 -3634 -1132
rect -3235 -1625 -3173 -882
rect -3235 -1693 -3173 -1687
rect -3278 -1834 -3216 -1822
rect -3294 -1916 -3284 -1834
rect -3204 -1916 -3194 -1834
rect -2466 -1844 -2420 -1220
rect -2336 -1720 -2092 -866
rect -2024 -1026 -2014 -970
rect -1956 -1026 -1946 -970
rect -2008 -1652 -1962 -1026
rect -1878 -1720 -1634 -866
rect -1550 -1844 -1504 -1220
rect -2484 -1904 -2474 -1844
rect -2412 -1904 -2402 -1844
rect -1568 -1904 -1558 -1844
rect -1496 -1904 -1486 -1844
rect -3746 -2356 -3736 -2264
rect -3640 -2356 -3630 -2264
rect -3794 -2533 -3744 -2388
rect -3955 -2643 -3744 -2533
rect -3955 -3190 -3845 -2643
rect -3794 -2788 -3744 -2643
rect -3714 -2818 -3668 -2356
rect -3636 -2558 -3584 -2388
rect -3278 -2558 -3216 -1916
rect -3100 -1958 -3035 -1952
rect -3100 -2160 -3035 -2023
rect -3107 -2166 -3029 -2160
rect -634 -2170 -588 -1222
rect -504 -1720 -260 -866
rect -176 -970 -130 -968
rect -192 -1026 -182 -970
rect -124 -1026 -114 -970
rect -176 -1662 -130 -1026
rect -46 -1720 198 -866
rect -2484 -2234 -2474 -2172
rect -2412 -2234 -2402 -2172
rect -1568 -2232 -1558 -2170
rect -1496 -2232 -1486 -2170
rect -652 -2232 -642 -2170
rect -580 -2232 -570 -2170
rect 282 -2174 328 -1214
rect 412 -1720 656 -866
rect 740 -970 786 -968
rect 724 -1026 734 -970
rect 792 -1026 802 -970
rect 740 -1662 786 -1026
rect 870 -1720 1114 -866
rect 1198 -2170 1244 -1212
rect 1328 -1720 1572 -866
rect 1656 -970 1702 -968
rect 1640 -1026 1650 -970
rect 1708 -1026 1718 -970
rect 1656 -1662 1702 -1026
rect 1786 -1720 2030 -866
rect 2090 -954 2166 8356
rect 2257 -664 2307 9744
rect 2416 1436 2472 9880
rect 2596 7486 2676 12436
rect 2783 8776 2833 12922
rect 9510 12582 9516 12642
rect 9576 12582 10826 12642
rect 3386 12446 3396 12498
rect 3520 12446 3530 12498
rect 3644 12446 3654 12498
rect 3778 12446 3788 12498
rect 3902 12446 3912 12498
rect 4036 12446 4046 12498
rect 4160 12446 4170 12498
rect 4294 12446 4304 12498
rect 4418 12446 4428 12498
rect 4552 12446 4562 12498
rect 4676 12446 4686 12498
rect 4810 12446 4820 12498
rect 4934 12446 4944 12498
rect 5068 12446 5078 12498
rect 5192 12446 5202 12498
rect 5326 12446 5336 12498
rect 5450 12446 5460 12498
rect 5584 12446 5594 12498
rect 5708 12446 5718 12498
rect 5842 12446 5852 12498
rect 5966 12446 5976 12498
rect 6100 12446 6110 12498
rect 6224 12446 6234 12498
rect 6358 12446 6368 12498
rect 6482 12446 6492 12498
rect 6616 12446 6626 12498
rect 6740 12446 6750 12498
rect 6874 12446 6884 12498
rect 6998 12446 7008 12498
rect 7132 12446 7142 12498
rect 7256 12446 7266 12498
rect 7390 12446 7400 12498
rect 7514 12446 7524 12498
rect 7648 12446 7658 12498
rect 7772 12446 7782 12498
rect 7906 12446 7916 12498
rect 8030 12446 8040 12498
rect 8164 12446 8174 12498
rect 8288 12446 8298 12498
rect 8422 12446 8432 12498
rect 3396 10524 3520 12446
rect 3560 10309 3614 12420
rect 3654 10524 3778 12446
rect 3822 12399 3868 12411
rect 3822 10623 3828 12399
rect 3862 10623 3868 12399
rect 3822 10611 3868 10623
rect 3912 10524 4036 12446
rect 3560 10249 3614 10255
rect 4076 10307 4130 12420
rect 4170 10524 4294 12446
rect 4428 10524 4552 12446
rect 4076 10247 4130 10253
rect 4592 10309 4646 12420
rect 4686 10524 4810 12446
rect 4854 12399 4900 12411
rect 4854 10623 4860 12399
rect 4894 10623 4900 12399
rect 4854 10611 4900 10623
rect 4944 10524 5068 12446
rect 4592 10249 4646 10255
rect 5108 10309 5162 12420
rect 5202 10524 5326 12446
rect 5460 10524 5584 12446
rect 5624 10439 5678 12420
rect 5718 10524 5842 12446
rect 5976 10524 6100 12446
rect 6140 10439 6194 12420
rect 6234 10524 6358 12446
rect 6492 10524 6616 12446
rect 5624 10385 6195 10439
rect 5108 10249 5162 10255
rect 3799 10201 3853 10207
rect 3550 9671 3600 9672
rect 3799 9671 3853 10147
rect 5883 10201 5937 10385
rect 6656 10307 6710 12420
rect 6750 10524 6874 12446
rect 6918 12399 6964 12411
rect 6918 10623 6924 12399
rect 6958 10623 6964 12399
rect 6918 10611 6964 10623
rect 7008 10524 7132 12446
rect 6656 10247 6710 10253
rect 6888 10310 6940 10316
rect 6888 10252 6940 10258
rect 7172 10309 7226 12420
rect 7266 10524 7390 12446
rect 7524 10524 7648 12446
rect 5883 10141 5937 10147
rect 6889 9673 6939 10252
rect 7172 10249 7226 10255
rect 7688 10309 7742 12420
rect 7782 10524 7906 12446
rect 7950 12399 7996 12411
rect 7950 10623 7956 12399
rect 7990 10623 7996 12399
rect 7950 10611 7996 10623
rect 8040 10524 8164 12446
rect 8204 10479 8258 12420
rect 8298 10524 8422 12446
rect 9596 10528 9640 12494
rect 9738 12448 9748 12500
rect 9800 12448 9810 12500
rect 9676 10606 9718 12418
rect 7688 10249 7742 10255
rect 8203 10392 8258 10479
rect 9678 10441 9716 10606
rect 9754 10528 9798 12448
rect 9838 10622 9872 12582
rect 9912 12500 9956 12502
rect 10070 12500 10114 12502
rect 9904 12448 9914 12500
rect 10112 12448 10122 12500
rect 9912 10528 9956 12448
rect 9994 10441 10032 12418
rect 10070 10528 10114 12448
rect 10154 10612 10188 12582
rect 10228 12500 10272 12502
rect 10386 12500 10430 12502
rect 10220 12448 10230 12500
rect 10428 12448 10438 12500
rect 10228 10528 10272 12448
rect 10310 10441 10348 12418
rect 10386 10528 10430 12448
rect 10470 10612 10504 12582
rect 10544 12500 10588 12502
rect 10702 12500 10746 12502
rect 10536 12448 10546 12500
rect 10744 12448 10754 12500
rect 10544 10528 10588 12448
rect 10626 10441 10664 12418
rect 10702 10528 10746 12448
rect 10786 10612 10820 12582
rect 10860 12500 10904 12502
rect 10852 12448 10862 12500
rect 10914 12448 10924 12500
rect 10860 10528 10904 12448
rect 10942 10441 10980 12418
rect 11018 10564 11060 12494
rect 11555 11546 11605 12922
rect 11808 12510 11880 12942
rect 12694 13018 12766 13024
rect 11808 12432 11880 12438
rect 12100 12105 12154 12688
rect 11825 12055 12154 12105
rect 11825 11556 11875 12055
rect 12100 11886 12154 12055
rect 12190 11850 12228 12760
rect 12266 12156 12320 12686
rect 12694 12274 12766 12946
rect 14149 12883 14159 12935
rect 14211 12883 14221 12935
rect 12926 12274 12972 12696
rect 12694 12202 12972 12274
rect 12266 12010 12308 12156
rect 12398 12124 12408 12156
rect 12398 12118 12412 12124
rect 12398 12040 12412 12046
rect 12398 12010 12408 12040
rect 12266 11884 12320 12010
rect 12926 11886 12972 12202
rect 12142 11768 12152 11850
rect 12260 11768 12270 11850
rect 13006 11848 13052 12764
rect 13086 11978 13132 12696
rect 13994 11978 14118 12644
rect 14160 12152 14210 12883
rect 14665 12882 14675 12934
rect 14727 12882 14737 12934
rect 14252 11978 14376 12644
rect 14510 11978 14634 12644
rect 14676 12151 14726 12882
rect 15697 12881 15707 12933
rect 15759 12881 15769 12933
rect 16213 12881 16223 12933
rect 16275 12881 16285 12933
rect 15181 12739 15191 12791
rect 15243 12739 15253 12791
rect 14768 11978 14892 12644
rect 15026 11978 15150 12644
rect 15192 12151 15242 12739
rect 15284 11978 15408 12644
rect 15542 11978 15666 12644
rect 15708 12151 15758 12881
rect 15800 11978 15924 12644
rect 16058 11978 16182 12644
rect 16224 12152 16274 12881
rect 16316 11978 16440 12644
rect 16971 12115 17037 13199
rect 17191 12929 17249 13341
rect 17191 12865 17249 12871
rect 16971 12043 17037 12049
rect 13086 11938 16440 11978
rect 13086 11886 13132 11938
rect 12966 11766 12976 11848
rect 13084 11766 13094 11848
rect 11548 11494 11554 11546
rect 11606 11494 11612 11546
rect 11800 11486 11810 11556
rect 11926 11486 11936 11556
rect 17467 11539 17529 13473
rect 20151 12943 20221 12949
rect 20151 12867 20221 12873
rect 18348 12801 18420 12807
rect 18098 12762 18148 12763
rect 18098 12729 18348 12762
rect 19904 12762 19954 12763
rect 20153 12762 20219 12867
rect 20935 12762 20985 12763
rect 18420 12729 18663 12762
rect 18098 12719 18663 12729
rect 18098 12138 18148 12719
rect 18190 12108 18314 12630
rect 18180 12056 18190 12108
rect 18314 12056 18324 12108
rect 18356 11969 18406 12549
rect 18448 12108 18572 12630
rect 18613 12137 18663 12719
rect 19388 12717 20985 12762
rect 18438 12056 18448 12108
rect 18572 12056 18582 12108
rect 18353 11906 18406 11969
rect 19130 11970 19180 12549
rect 19222 12108 19346 12630
rect 19388 12137 19438 12717
rect 19480 12108 19604 12630
rect 19212 12056 19222 12108
rect 19346 12056 19356 12108
rect 19470 12056 19480 12108
rect 19604 12056 19614 12108
rect 19646 11970 19696 12549
rect 19738 12108 19862 12630
rect 19904 12138 19954 12717
rect 19996 12108 20120 12630
rect 19728 12056 19738 12108
rect 19862 12056 19872 12108
rect 19986 12056 19996 12108
rect 20120 12056 20130 12108
rect 20162 11970 20212 12549
rect 20254 12108 20378 12630
rect 20420 12137 20470 12717
rect 20512 12108 20636 12630
rect 20244 12056 20254 12108
rect 20378 12056 20388 12108
rect 20502 12056 20512 12108
rect 20636 12056 20646 12108
rect 20678 11970 20728 12549
rect 20770 12108 20894 12630
rect 20935 12138 20985 12717
rect 21028 12108 21152 12630
rect 20760 12056 20770 12108
rect 20894 12056 20904 12108
rect 21018 12056 21028 12108
rect 21152 12056 21162 12108
rect 21194 11970 21244 12549
rect 22970 12543 23094 12630
rect 22727 12231 23094 12543
rect 22200 12225 22279 12231
rect 19130 11968 22091 11970
rect 19130 11924 22105 11968
rect 18353 11552 18403 11906
rect 22032 11878 22105 11924
rect 22030 11846 22105 11878
rect 18352 11546 18404 11552
rect 18352 11488 18404 11494
rect 17467 11471 17529 11477
rect 11684 11400 11756 11406
rect 19953 11367 20016 11373
rect 11550 11230 11622 11236
rect 8203 10309 8257 10392
rect 9666 10379 10985 10441
rect 8203 10249 8257 10255
rect 9770 9932 9822 9938
rect 9770 9874 9822 9880
rect 9554 9802 9606 9808
rect 9554 9744 9606 9750
rect 4066 9671 4116 9672
rect 3549 9621 4116 9671
rect 5097 9623 8760 9673
rect 3374 9486 3384 9538
rect 3508 9486 3518 9538
rect 2780 8432 2856 8776
rect 2780 8350 2856 8356
rect 2596 7480 2688 7486
rect 2596 7428 2636 7480
rect 3292 7483 3342 9460
rect 3384 7564 3508 9486
rect 3550 7644 3600 9621
rect 3799 9619 3853 9621
rect 3632 9486 3642 9538
rect 3766 9486 3776 9538
rect 3890 9486 3900 9538
rect 4024 9486 4034 9538
rect 3642 7564 3766 9486
rect 3808 7486 3858 9460
rect 3900 7564 4024 9486
rect 4066 7644 4116 9621
rect 4148 9486 4158 9538
rect 4282 9486 4292 9538
rect 4922 9486 4932 9538
rect 5056 9486 5066 9538
rect 4158 7564 4282 9486
rect 3808 7483 3864 7486
rect 4324 7483 4374 9460
rect 3292 7480 4375 7483
rect 3292 7433 3812 7480
rect 3292 7432 3342 7433
rect 3808 7432 3812 7433
rect 2596 7422 2688 7428
rect 3864 7433 4375 7480
rect 4840 7480 4890 9460
rect 4932 7564 5056 9486
rect 5098 7644 5148 9623
rect 5180 9486 5190 9538
rect 5314 9486 5324 9538
rect 5438 9486 5448 9538
rect 5572 9486 5582 9538
rect 5190 7564 5314 9486
rect 5356 7480 5406 9460
rect 5448 7564 5572 9486
rect 5614 7644 5664 9623
rect 5696 9486 5706 9538
rect 5830 9486 5840 9538
rect 5954 9486 5964 9538
rect 6088 9486 6098 9538
rect 5706 7564 5830 9486
rect 5872 7480 5922 9460
rect 5964 7564 6088 9486
rect 6130 7644 6180 9623
rect 6212 9486 6222 9538
rect 6346 9486 6356 9538
rect 6470 9486 6480 9538
rect 6604 9486 6614 9538
rect 6222 7564 6346 9486
rect 6388 7480 6438 9460
rect 6480 7564 6604 9486
rect 6646 7644 6696 9623
rect 6728 9486 6738 9538
rect 6862 9486 6872 9538
rect 6986 9486 6996 9538
rect 7120 9486 7130 9538
rect 6738 7564 6862 9486
rect 6602 7504 6718 7510
rect 6484 7480 6602 7504
rect 4324 7432 4374 7433
rect 4840 7432 6602 7480
rect 4840 7431 4890 7432
rect 3812 7422 3864 7428
rect 2596 7368 2687 7422
rect 6484 7388 6602 7432
rect 6904 7480 6954 9460
rect 6996 7564 7120 9486
rect 7162 7644 7212 9623
rect 7244 9486 7254 9538
rect 7378 9486 7388 9538
rect 7502 9486 7512 9538
rect 7636 9486 7646 9538
rect 7254 7564 7378 9486
rect 7420 7480 7470 9460
rect 7512 7564 7636 9486
rect 7678 7644 7728 9623
rect 7760 9486 7770 9538
rect 7894 9486 7904 9538
rect 8018 9486 8028 9538
rect 8152 9486 8162 9538
rect 7770 7564 7894 9486
rect 7936 7480 7986 9460
rect 8028 7564 8152 9486
rect 8194 7644 8244 9623
rect 8276 9486 8286 9538
rect 8410 9486 8420 9538
rect 8534 9486 8544 9538
rect 8668 9486 8678 9538
rect 8286 7564 8410 9486
rect 8452 7480 8502 9460
rect 8544 7564 8668 9486
rect 8710 7644 8760 9623
rect 8792 9486 8802 9538
rect 8926 9486 8936 9538
rect 8802 7564 8926 9486
rect 8968 7480 9018 9460
rect 9555 8422 9605 9744
rect 9554 8416 9606 8422
rect 9554 8358 9606 8364
rect 9771 8280 9821 9874
rect 9770 8274 9822 8280
rect 9770 8216 9822 8222
rect 6718 7432 9020 7480
rect 10213 7463 10275 10379
rect 10213 7395 10275 7401
rect 10898 8591 10977 8597
rect 6602 7382 6718 7388
rect 2637 5876 2687 7368
rect 10280 7210 10344 7216
rect 10138 6954 10190 6960
rect 3336 6778 9958 6830
rect 2608 5792 2618 5876
rect 2698 5792 2708 5876
rect 2637 1584 2687 5792
rect 3244 5394 3254 6616
rect 3310 5394 3320 6616
rect 3348 5320 3474 6778
rect 3502 5394 3512 6616
rect 3568 5394 3578 6616
rect 3606 5320 3732 6778
rect 3760 5394 3770 6616
rect 3826 5394 3836 6616
rect 3864 5230 3990 6696
rect 4018 5394 4028 6616
rect 4084 5394 4094 6616
rect 4122 5230 4248 6696
rect 4276 5394 4286 6616
rect 4342 5394 4352 6616
rect 4380 5230 4506 6696
rect 4534 5394 4544 6616
rect 4600 5394 4610 6616
rect 4638 5230 4764 6696
rect 4792 5394 4802 6616
rect 4858 5394 4868 6616
rect 4896 5320 5022 6778
rect 5050 5394 5060 6616
rect 5116 5394 5126 6616
rect 5154 5320 5280 6778
rect 5308 5394 5318 6616
rect 5374 5394 5384 6616
rect 5412 5320 5538 6778
rect 5566 5394 5576 6616
rect 5632 5394 5642 6616
rect 5670 5320 5796 6778
rect 5824 5394 5834 6616
rect 5890 5394 5900 6616
rect 5928 5230 6054 6696
rect 6082 5394 6092 6616
rect 6148 5394 6158 6616
rect 6186 5230 6312 6696
rect 6340 5394 6350 6616
rect 6406 5394 6416 6616
rect 6444 5230 6570 6696
rect 6598 5394 6608 6616
rect 6664 5394 6674 6616
rect 6702 5230 6828 6696
rect 6856 5394 6866 6616
rect 6922 5394 6932 6616
rect 6960 5320 7086 6778
rect 7114 5394 7124 6616
rect 7180 5394 7190 6616
rect 7218 5320 7344 6778
rect 7372 5394 7382 6616
rect 7438 5394 7448 6616
rect 7476 5320 7602 6778
rect 7630 5394 7640 6616
rect 7696 5394 7706 6616
rect 7734 5320 7860 6778
rect 7888 5394 7898 6616
rect 7954 5394 7964 6616
rect 7992 5230 8118 6696
rect 8146 5394 8156 6616
rect 8212 5394 8222 6616
rect 8250 5230 8376 6696
rect 8404 5394 8414 6616
rect 8470 5394 8480 6616
rect 8508 5230 8634 6696
rect 8662 5394 8672 6616
rect 8728 5394 8738 6616
rect 8766 5230 8892 6696
rect 8920 5394 8930 6616
rect 8986 5394 8996 6616
rect 9024 5320 9150 6778
rect 9178 5394 9188 6616
rect 9244 5394 9254 6616
rect 9282 5320 9408 6778
rect 9436 5394 9446 6616
rect 9502 5394 9512 6616
rect 2836 5182 9740 5230
rect 2836 3062 2884 5182
rect 3244 3790 3254 5012
rect 3310 3790 3320 5012
rect 3348 3716 3474 5182
rect 3502 3790 3512 5012
rect 3568 3790 3578 5012
rect 3606 3716 3732 5182
rect 3760 3790 3770 5012
rect 3826 3790 3836 5012
rect 3864 3628 3990 5092
rect 4018 3790 4028 5012
rect 4084 3790 4094 5012
rect 4122 3628 4248 5092
rect 4276 3790 4286 5012
rect 4342 3790 4352 5012
rect 4380 3628 4506 5092
rect 4534 3790 4544 5012
rect 4600 3790 4610 5012
rect 4638 3628 4764 5092
rect 4792 3790 4802 5012
rect 4858 3790 4868 5012
rect 4896 3716 5022 5182
rect 5050 3790 5060 5012
rect 5116 3790 5126 5012
rect 5154 3716 5280 5182
rect 5308 3790 5318 5012
rect 5374 3790 5384 5012
rect 5412 3716 5538 5182
rect 5566 3790 5576 5012
rect 5632 3790 5642 5012
rect 5670 3716 5796 5182
rect 5824 3790 5834 5012
rect 5890 3790 5900 5012
rect 5928 3628 6054 5092
rect 6082 3790 6092 5012
rect 6148 3790 6158 5012
rect 6186 3628 6312 5092
rect 6340 3790 6350 5012
rect 6406 3790 6416 5012
rect 6444 3628 6570 5092
rect 6598 3790 6608 5012
rect 6664 3790 6674 5012
rect 6702 3628 6828 5092
rect 6856 3790 6866 5012
rect 6922 3790 6932 5012
rect 6960 3716 7086 5182
rect 7114 3790 7124 5012
rect 7180 3790 7190 5012
rect 7218 3716 7344 5182
rect 7372 3790 7382 5012
rect 7438 3790 7448 5012
rect 7476 3716 7602 5182
rect 7630 3790 7640 5012
rect 7696 3790 7706 5012
rect 7734 3716 7860 5182
rect 7888 3790 7898 5012
rect 7954 3790 7964 5012
rect 7992 3628 8118 5092
rect 8146 3790 8156 5012
rect 8212 3790 8222 5012
rect 8250 3628 8376 5092
rect 8404 3790 8414 5012
rect 8470 3790 8480 5012
rect 8508 3628 8634 5092
rect 8662 3790 8672 5012
rect 8728 3790 8738 5012
rect 8766 3628 8892 5092
rect 8920 3790 8930 5012
rect 8986 3790 8996 5012
rect 9024 3716 9150 5182
rect 9178 3790 9188 5012
rect 9244 3790 9254 5012
rect 9282 3716 9408 5182
rect 9436 3790 9446 5012
rect 9502 3790 9512 5012
rect 9906 3648 9958 6778
rect 3346 3626 9426 3628
rect 9906 3626 9980 3648
rect 3346 3576 9980 3626
rect 9348 3574 9980 3576
rect 6035 3346 6041 3425
rect 6120 3346 6126 3425
rect 2834 3056 2886 3062
rect 2834 2998 2886 3004
rect 4760 1946 4812 1952
rect 4760 1888 4812 1894
rect 3450 1826 3522 1832
rect 2636 1578 2688 1584
rect 2636 1520 2688 1526
rect 2416 1374 2472 1380
rect 3450 880 3522 1754
rect 2840 838 4138 880
rect 2756 -316 2800 732
rect 2840 -246 2874 838
rect 2914 -296 2958 740
rect 2892 -348 2902 -296
rect 2958 -348 2968 -296
rect 2998 -418 3032 662
rect 3072 -296 3116 740
rect 3156 -246 3190 838
rect 3450 836 3522 838
rect 3230 -296 3274 740
rect 3062 -348 3072 -296
rect 3274 -348 3284 -296
rect 3136 -414 3220 -408
rect 3094 -418 3100 -414
rect 2998 -464 3100 -418
rect 3094 -466 3100 -464
rect 3314 -418 3348 662
rect 3388 -296 3432 740
rect 3472 -246 3506 836
rect 3546 -296 3590 740
rect 3378 -348 3388 -296
rect 3590 -348 3600 -296
rect 3630 -418 3664 662
rect 3704 -296 3748 740
rect 3788 -246 3822 838
rect 3862 -296 3906 740
rect 3694 -348 3704 -296
rect 3906 -348 3916 -296
rect 3946 -418 3980 662
rect 4020 -296 4064 740
rect 4104 -246 4138 838
rect 4010 -348 4020 -296
rect 4076 -348 4086 -296
rect 4178 -316 4222 740
rect 4762 -280 4810 1888
rect 5518 1578 5570 1584
rect 5518 1520 5570 1526
rect 5378 1436 5434 1442
rect 4905 1186 5007 1187
rect 4888 876 4898 1186
rect 5010 876 5020 1186
rect 4748 -286 4820 -280
rect 3220 -464 3882 -418
rect 3136 -472 3220 -466
rect 3872 -476 3882 -464
rect 4004 -476 4014 -418
rect 2256 -670 2308 -664
rect 2256 -728 2308 -722
rect 2234 -866 2244 -812
rect 2488 -866 2498 -812
rect 2692 -866 2702 -812
rect 2946 -866 2956 -812
rect 3150 -866 3160 -812
rect 3404 -866 3414 -812
rect 3608 -866 3618 -812
rect 3862 -866 3872 -812
rect 2082 -960 2172 -954
rect 2082 -1036 2090 -960
rect 2166 -1036 2172 -960
rect 2082 -1044 2172 -1036
rect -3107 -2250 -3029 -2244
rect -3636 -2624 -3216 -2558
rect -3636 -2786 -3584 -2624
rect -3748 -2910 -3738 -2818
rect -3642 -2910 -3632 -2818
rect -3278 -3038 -3216 -2624
rect -2466 -2848 -2420 -2234
rect -3292 -3120 -3282 -3038
rect -3202 -3120 -3192 -3038
rect -2280 -3204 -2150 -2350
rect -2280 -3290 -2264 -3204
rect -2170 -3290 -2150 -3204
rect -1820 -3204 -1690 -2350
rect -1550 -2848 -1504 -2232
rect -1820 -3290 -1804 -3204
rect -1710 -3290 -1690 -3204
rect -1358 -3202 -1228 -2348
rect -1358 -3288 -1340 -3202
rect -1246 -3288 -1228 -3202
rect -902 -3194 -772 -2340
rect -634 -2848 -588 -2232
rect 246 -2242 256 -2174
rect 352 -2242 362 -2174
rect 1180 -2232 1190 -2170
rect 1252 -2232 1262 -2170
rect 2114 -2176 2160 -1214
rect 2244 -1720 2488 -866
rect 2572 -970 2618 -968
rect 2556 -1026 2566 -970
rect 2624 -1026 2634 -970
rect 2572 -1662 2618 -1026
rect 2702 -1720 2946 -866
rect -902 -3280 -886 -3194
rect -792 -3280 -772 -3194
rect -450 -3204 -320 -2350
rect -450 -3290 -432 -3204
rect -338 -3290 -320 -3204
rect 14 -3204 144 -2350
rect 282 -2958 328 -2436
rect 260 -2962 348 -2958
rect 250 -3108 260 -2962
rect 348 -3108 358 -2962
rect 270 -3112 338 -3108
rect 14 -3290 30 -3204
rect 124 -3290 144 -3204
rect 466 -3206 596 -2352
rect 466 -3292 482 -3206
rect 576 -3292 596 -3206
rect 930 -3204 1060 -2352
rect 1198 -2848 1244 -2232
rect 2096 -2238 2106 -2176
rect 2168 -2238 2178 -2176
rect 3030 -2178 3076 -1214
rect 3160 -1720 3404 -866
rect 3488 -970 3534 -968
rect 3472 -1026 3482 -970
rect 3540 -1026 3550 -970
rect 3488 -1662 3534 -1026
rect 3618 -1720 3862 -866
rect 4748 -1054 4820 -358
rect 4918 -408 4994 876
rect 5378 106 5434 1380
rect 5519 172 5569 1520
rect 6041 1471 6120 3346
rect 9928 2898 9980 3574
rect 10138 3534 10190 6902
rect 10280 4988 10344 7146
rect 10898 7051 10977 8512
rect 10898 6997 10915 7051
rect 10969 6997 10977 7051
rect 10449 5234 10507 5240
rect 10274 4982 10350 4988
rect 10274 4918 10280 4982
rect 10344 4918 10350 4982
rect 10274 4910 10350 4918
rect 10138 3476 10190 3482
rect 10449 3535 10507 5176
rect 10449 3471 10507 3477
rect 10898 3425 10977 6997
rect 11184 8082 11256 8088
rect 11034 6956 11086 6962
rect 11034 5118 11086 6904
rect 11184 5288 11256 8010
rect 11550 8082 11622 11158
rect 11684 9548 11756 11328
rect 11684 9470 11756 9476
rect 12222 11351 12272 11352
rect 12738 11351 12788 11352
rect 13770 11351 13820 11352
rect 15318 11351 15368 11352
rect 15834 11351 15884 11352
rect 17898 11351 17948 11352
rect 18414 11351 18464 11352
rect 12222 11304 19953 11351
rect 20994 11351 21044 11352
rect 21510 11351 21560 11352
rect 20016 11304 21561 11351
rect 12222 11301 21561 11304
rect 12222 8726 12272 11301
rect 12304 11168 12314 11220
rect 12438 11168 12448 11220
rect 12562 11168 12572 11220
rect 12696 11168 12706 11220
rect 12314 8646 12438 11168
rect 12572 8646 12696 11168
rect 12738 8726 12788 11301
rect 12820 11168 12830 11220
rect 12954 11168 12964 11220
rect 13078 11168 13088 11220
rect 13212 11168 13222 11220
rect 13336 11168 13346 11220
rect 13470 11168 13480 11220
rect 13594 11168 13604 11220
rect 13728 11168 13738 11220
rect 12830 8646 12954 11168
rect 12998 11121 13044 11133
rect 12998 8745 13004 11121
rect 13038 8745 13044 11121
rect 12998 8733 13044 8745
rect 13088 8646 13212 11168
rect 13254 8583 13304 11140
rect 13346 8646 13470 11168
rect 13514 11121 13560 11133
rect 13514 8745 13520 11121
rect 13554 8745 13560 11121
rect 13514 8733 13560 8745
rect 13604 8646 13728 11168
rect 13770 8726 13820 11301
rect 13852 11168 13862 11220
rect 13986 11168 13996 11220
rect 14110 11168 14120 11220
rect 14244 11168 14254 11220
rect 14368 11168 14378 11220
rect 14502 11168 14512 11220
rect 14626 11168 14636 11220
rect 14760 11168 14770 11220
rect 14884 11168 14894 11220
rect 15018 11168 15028 11220
rect 15142 11168 15152 11220
rect 15276 11168 15286 11220
rect 13862 8646 13986 11168
rect 14030 11121 14076 11133
rect 14030 8745 14036 11121
rect 14070 8745 14076 11121
rect 14030 8733 14076 8745
rect 14120 8646 14244 11168
rect 13666 8591 13745 8597
rect 13254 8533 13666 8583
rect 13254 8532 13304 8533
rect 14286 8583 14336 11140
rect 14378 8646 14502 11168
rect 14546 11121 14592 11133
rect 14546 8745 14552 11121
rect 14586 8745 14592 11121
rect 14546 8733 14592 8745
rect 14636 8646 14760 11168
rect 14802 8583 14852 11140
rect 14894 8646 15018 11168
rect 15062 11121 15108 11133
rect 15062 8745 15068 11121
rect 15102 8745 15108 11121
rect 15062 8733 15108 8745
rect 15152 8646 15276 11168
rect 15318 8726 15368 11301
rect 15400 11168 15410 11220
rect 15534 11168 15544 11220
rect 15658 11168 15668 11220
rect 15792 11168 15802 11220
rect 15410 8646 15534 11168
rect 15668 8646 15792 11168
rect 15834 8726 15884 11301
rect 15916 11168 15926 11220
rect 16050 11168 16060 11220
rect 16174 11168 16184 11220
rect 16308 11168 16318 11220
rect 16432 11168 16442 11220
rect 16566 11168 16576 11220
rect 16690 11168 16700 11220
rect 16824 11168 16834 11220
rect 16948 11168 16958 11220
rect 17082 11168 17092 11220
rect 17206 11168 17216 11220
rect 17340 11168 17350 11220
rect 17464 11168 17474 11220
rect 17598 11168 17608 11220
rect 17722 11168 17732 11220
rect 17856 11168 17866 11220
rect 15926 8646 16050 11168
rect 16094 11121 16140 11133
rect 16094 8745 16100 11121
rect 16134 8745 16140 11121
rect 16094 8733 16140 8745
rect 16184 8646 16308 11168
rect 16350 8583 16400 11140
rect 16442 8646 16566 11168
rect 16610 11121 16656 11133
rect 16610 8745 16616 11121
rect 16650 8745 16656 11121
rect 16610 8733 16656 8745
rect 16700 8646 16824 11168
rect 16866 8583 16916 11140
rect 16958 8646 17082 11168
rect 17126 11121 17172 11133
rect 17126 8745 17132 11121
rect 17166 8745 17172 11121
rect 17126 8733 17172 8745
rect 17216 8646 17340 11168
rect 17382 8583 17432 11140
rect 17474 8646 17598 11168
rect 17642 11121 17688 11133
rect 17642 8745 17648 11121
rect 17682 8745 17688 11121
rect 17642 8733 17688 8745
rect 17732 8646 17856 11168
rect 17898 8726 17948 11301
rect 17980 11168 17990 11220
rect 18114 11168 18124 11220
rect 18238 11168 18248 11220
rect 18372 11168 18382 11220
rect 17990 8646 18114 11168
rect 18248 8646 18372 11168
rect 18414 8726 18464 11301
rect 19953 11298 20016 11301
rect 18496 11168 18506 11220
rect 18630 11168 18640 11220
rect 18754 11168 18764 11220
rect 18888 11168 18898 11220
rect 19012 11168 19022 11220
rect 19146 11168 19156 11220
rect 19270 11168 19280 11220
rect 19404 11168 19414 11220
rect 19528 11168 19538 11220
rect 19662 11168 19672 11220
rect 19786 11168 19796 11220
rect 19920 11168 19930 11220
rect 18506 8646 18630 11168
rect 18674 11121 18720 11133
rect 18674 8745 18680 11121
rect 18714 8745 18720 11121
rect 18674 8733 18720 8745
rect 18764 8646 18888 11168
rect 18930 8583 18980 11140
rect 19022 8646 19146 11168
rect 19190 11121 19236 11133
rect 19190 8745 19196 11121
rect 19230 8745 19236 11121
rect 19190 8733 19236 8745
rect 19280 8646 19404 11168
rect 19446 8583 19496 11140
rect 19538 8646 19662 11168
rect 19706 11121 19752 11133
rect 19706 8745 19712 11121
rect 19746 8745 19752 11121
rect 19706 8733 19752 8745
rect 19796 8646 19920 11168
rect 19962 8726 20012 11298
rect 20044 11168 20054 11220
rect 20178 11168 20188 11220
rect 20302 11168 20312 11220
rect 20436 11168 20446 11220
rect 20560 11168 20570 11220
rect 20694 11168 20704 11220
rect 20818 11168 20828 11220
rect 20952 11168 20962 11220
rect 20054 8646 20178 11168
rect 20222 11121 20268 11133
rect 20222 8745 20228 11121
rect 20262 8745 20268 11121
rect 20222 8733 20268 8745
rect 20312 8646 20436 11168
rect 20478 8583 20528 11140
rect 20570 8646 20694 11168
rect 20738 11121 20784 11133
rect 20738 8745 20744 11121
rect 20778 8745 20784 11121
rect 20738 8733 20784 8745
rect 20828 8646 20952 11168
rect 20994 8726 21044 11301
rect 21076 11168 21086 11220
rect 21210 11168 21220 11220
rect 21334 11168 21344 11220
rect 21468 11168 21478 11220
rect 21086 8646 21210 11168
rect 21344 8646 21468 11168
rect 21510 8726 21560 11301
rect 13745 8533 20529 8583
rect 14286 8532 14336 8533
rect 14802 8532 14852 8533
rect 16350 8532 16400 8533
rect 16866 8532 16916 8533
rect 17382 8532 17432 8533
rect 18930 8532 18980 8533
rect 19446 8532 19496 8533
rect 20478 8532 20528 8533
rect 13666 8506 13745 8512
rect 13672 8074 13733 8506
rect 18683 8160 18746 8166
rect 11974 8011 16161 8074
rect 18683 8072 18746 8097
rect 11550 8004 11622 8010
rect 11804 7886 11814 7938
rect 11938 7886 11948 7938
rect 11722 5281 11772 7858
rect 11814 5364 11938 7886
rect 11980 5444 12030 8011
rect 12062 7886 12072 7938
rect 12196 7886 12206 7938
rect 12320 7886 12330 7938
rect 12454 7886 12464 7938
rect 12072 5364 12196 7886
rect 12236 5281 12286 7858
rect 12330 5364 12454 7886
rect 12496 5444 12546 8011
rect 12578 7886 12588 7938
rect 12712 7886 12722 7938
rect 12836 7886 12846 7938
rect 12970 7886 12980 7938
rect 12588 5364 12712 7886
rect 12754 5281 12804 7858
rect 12846 5364 12970 7886
rect 13012 5444 13062 8011
rect 13094 7886 13104 7938
rect 13228 7886 13238 7938
rect 13352 7886 13362 7938
rect 13486 7886 13496 7938
rect 13104 5364 13228 7886
rect 13268 5282 13318 7858
rect 13362 5364 13486 7886
rect 13528 5444 13578 8011
rect 13610 7886 13620 7938
rect 13744 7886 13754 7938
rect 13868 7886 13878 7938
rect 14002 7886 14012 7938
rect 13620 5364 13744 7886
rect 13268 5281 13368 5282
rect 13786 5281 13836 7858
rect 13878 5364 14002 7886
rect 14044 5444 14094 8011
rect 14126 7886 14136 7938
rect 14260 7886 14270 7938
rect 14384 7886 14394 7938
rect 14518 7886 14528 7938
rect 14136 5364 14260 7886
rect 14300 5294 14350 7858
rect 14394 5364 14518 7886
rect 14560 5444 14610 8011
rect 14642 7886 14652 7938
rect 14776 7886 14786 7938
rect 14900 7886 14910 7938
rect 15034 7886 15044 7938
rect 14652 5364 14776 7886
rect 14288 5288 14360 5294
rect 11721 5231 14288 5281
rect 11184 5210 11256 5216
rect 11034 5060 11086 5066
rect 10898 3340 10977 3346
rect 6041 1386 6120 1392
rect 6287 2553 6357 2559
rect 6287 352 6357 2483
rect 9928 2442 9980 2846
rect 11195 2703 11253 5210
rect 13144 5120 13199 5126
rect 12759 4991 12829 4997
rect 12560 4816 12612 4822
rect 12560 4758 12612 4764
rect 12415 4585 12481 4591
rect 12415 2797 12481 4519
rect 12562 3168 12610 4758
rect 12560 3162 12612 3168
rect 12560 3104 12612 3110
rect 12415 2725 12481 2731
rect 11195 2639 11253 2645
rect 12759 2564 12829 4921
rect 12994 3534 13046 3540
rect 12994 2822 13046 3482
rect 12994 2764 13046 2770
rect 13144 2686 13199 5065
rect 13316 3384 13368 5231
rect 14818 5281 14868 7858
rect 14910 5364 15034 7886
rect 15076 5444 15126 8011
rect 15158 7886 15168 7938
rect 15292 7886 15302 7938
rect 15416 7886 15426 7938
rect 15550 7886 15560 7938
rect 15168 5364 15292 7886
rect 15332 5281 15384 7858
rect 15426 5364 15550 7886
rect 15592 5444 15642 8011
rect 15674 7886 15684 7938
rect 15808 7886 15818 7938
rect 15932 7886 15942 7938
rect 16066 7886 16076 7938
rect 15684 5364 15808 7886
rect 15848 5281 15900 7858
rect 15942 5364 16066 7886
rect 16108 5444 16158 8011
rect 17134 8009 21326 8072
rect 16190 7886 16200 7938
rect 16324 7886 16334 7938
rect 16964 7886 16974 7938
rect 17098 7886 17108 7938
rect 16200 5364 16324 7886
rect 16366 5281 16416 7858
rect 16882 5281 16932 7858
rect 16974 5364 17098 7886
rect 17140 5444 17190 8009
rect 17222 7886 17232 7938
rect 17356 7886 17366 7938
rect 17480 7886 17490 7938
rect 17614 7886 17624 7938
rect 17232 5364 17356 7886
rect 17396 5281 17446 7858
rect 17490 5364 17614 7886
rect 17656 5444 17706 8009
rect 17738 7886 17748 7938
rect 17872 7886 17882 7938
rect 17996 7886 18006 7938
rect 18130 7886 18140 7938
rect 17748 5364 17872 7886
rect 17914 5281 17964 7858
rect 18006 5364 18130 7886
rect 18172 5444 18222 8009
rect 18254 7886 18264 7938
rect 18388 7886 18398 7938
rect 18512 7886 18522 7938
rect 18646 7886 18656 7938
rect 18264 5364 18388 7886
rect 18428 5281 18478 7858
rect 18522 5364 18646 7886
rect 18688 5444 18738 8009
rect 18770 7886 18780 7938
rect 18904 7886 18914 7938
rect 19028 7886 19038 7938
rect 19162 7886 19172 7938
rect 18780 5364 18904 7886
rect 18946 5281 18996 7858
rect 19038 5364 19162 7886
rect 19204 5444 19254 8009
rect 19286 7886 19296 7938
rect 19420 7886 19430 7938
rect 19544 7886 19554 7938
rect 19678 7886 19688 7938
rect 19296 5364 19420 7886
rect 19460 5281 19510 7858
rect 19554 5364 19678 7886
rect 19720 5444 19770 8009
rect 19802 7886 19812 7938
rect 19936 7886 19946 7938
rect 20060 7886 20070 7938
rect 20194 7886 20204 7938
rect 19812 5364 19936 7886
rect 19978 5281 20028 7858
rect 20070 5364 20194 7886
rect 20236 5444 20286 8009
rect 20318 7886 20328 7938
rect 20452 7886 20462 7938
rect 20576 7886 20586 7938
rect 20710 7886 20720 7938
rect 20328 5364 20452 7886
rect 20492 5281 20544 7858
rect 20586 5364 20710 7886
rect 20752 5444 20802 8009
rect 20834 7886 20844 7938
rect 20968 7886 20978 7938
rect 21092 7886 21102 7938
rect 21226 7886 21236 7938
rect 20844 5364 20968 7886
rect 21008 5281 21060 7858
rect 21102 5364 21226 7886
rect 21268 5444 21318 8009
rect 21350 7886 21360 7938
rect 21484 7886 21494 7938
rect 21360 5364 21484 7886
rect 21526 5281 21576 7858
rect 14360 5231 16416 5281
rect 16881 5231 21576 5281
rect 14288 5210 14360 5216
rect 13880 4709 13930 4710
rect 14396 4709 14446 4710
rect 14645 4709 14695 5231
rect 16192 4824 16244 4830
rect 16192 4766 16244 4772
rect 17270 4828 17322 4834
rect 19201 4830 19251 5231
rect 17270 4770 17322 4776
rect 19200 4824 19252 4830
rect 14912 4709 14962 4710
rect 15428 4709 15478 4710
rect 13880 4659 15478 4709
rect 13880 3646 13930 4659
rect 13962 4526 13972 4578
rect 14096 4526 14106 4578
rect 14220 4526 14230 4578
rect 14354 4526 14364 4578
rect 13972 3564 14096 4526
rect 14138 3483 14188 4496
rect 14230 3564 14354 4526
rect 14396 3646 14446 4659
rect 14478 4526 14488 4578
rect 14612 4526 14622 4578
rect 14736 4526 14746 4578
rect 14870 4526 14880 4578
rect 14488 3564 14612 4526
rect 14654 3483 14704 4496
rect 14746 3564 14870 4526
rect 14912 3646 14962 4659
rect 14994 4526 15004 4578
rect 15128 4526 15138 4578
rect 15252 4526 15262 4578
rect 15386 4526 15396 4578
rect 15004 3564 15128 4526
rect 15170 3483 15220 4496
rect 15262 3564 15386 4526
rect 15428 3646 15478 4659
rect 15944 4709 15994 4710
rect 16193 4709 16243 4766
rect 15944 4708 16509 4709
rect 15944 4659 16510 4708
rect 15944 3646 15994 4659
rect 16193 4655 16243 4659
rect 16026 4526 16036 4578
rect 16160 4526 16170 4578
rect 16284 4526 16294 4578
rect 16418 4526 16428 4578
rect 16036 3564 16160 4526
rect 14138 3433 15220 3483
rect 14138 3432 14188 3433
rect 14654 3432 14751 3433
rect 15170 3432 15220 3433
rect 16202 3483 16252 4496
rect 16294 3564 16418 4526
rect 16460 3644 16510 4659
rect 16542 4526 16552 4578
rect 16676 4526 16686 4578
rect 16552 3564 16676 4526
rect 16718 3483 16768 4496
rect 16202 3433 16768 3483
rect 16202 3432 16252 3433
rect 13316 3326 13368 3332
rect 13144 2625 13199 2631
rect 13660 2822 13712 2828
rect 12759 2488 12829 2494
rect 12914 2442 13542 2454
rect 6904 2390 13542 2442
rect 6820 1618 6830 2230
rect 6884 1618 6894 2230
rect 6924 1546 7048 2390
rect 7078 1618 7088 2230
rect 7142 1618 7152 2230
rect 7182 1546 7306 2390
rect 7336 1618 7346 2230
rect 7400 1618 7410 2230
rect 7440 1454 7564 2302
rect 7594 1618 7604 2230
rect 7658 1618 7668 2230
rect 7698 1454 7822 2302
rect 7852 1618 7862 2230
rect 7916 1618 7926 2230
rect 7956 1454 8080 2302
rect 8110 1618 8120 2230
rect 8174 1618 8184 2230
rect 8214 1454 8338 2302
rect 8368 1618 8378 2230
rect 8432 1618 8442 2230
rect 8472 1546 8596 2390
rect 8626 1618 8636 2230
rect 8690 1618 8700 2230
rect 8730 1546 8854 2390
rect 8884 1618 8894 2230
rect 8948 1618 8958 2230
rect 8988 1546 9112 2390
rect 9142 1618 9152 2230
rect 9206 1618 9216 2230
rect 9246 1546 9370 2390
rect 9400 1618 9410 2230
rect 9464 1618 9474 2230
rect 9504 1454 9628 2302
rect 9658 1618 9668 2230
rect 9722 1618 9732 2230
rect 9762 1454 9886 2302
rect 9916 1618 9926 2230
rect 9980 1618 9990 2230
rect 10020 1454 10144 2302
rect 10174 1618 10184 2230
rect 10238 1618 10248 2230
rect 10278 1454 10402 2302
rect 10432 1618 10442 2230
rect 10496 1618 10506 2230
rect 10536 1546 10660 2390
rect 10690 1618 10700 2230
rect 10754 1618 10764 2230
rect 10794 1546 10918 2390
rect 10948 1618 10958 2230
rect 11012 1618 11022 2230
rect 11052 1546 11176 2390
rect 11206 1618 11216 2230
rect 11270 1618 11280 2230
rect 11310 1546 11434 2390
rect 11464 1618 11474 2230
rect 11528 1618 11538 2230
rect 11568 1454 11692 2302
rect 11722 1618 11732 2230
rect 11786 1618 11796 2230
rect 11826 1454 11950 2302
rect 11980 1618 11990 2230
rect 12044 1618 12054 2230
rect 12084 1454 12208 2302
rect 12238 1618 12248 2230
rect 12302 1618 12312 2230
rect 12342 1454 12466 2302
rect 12496 1618 12506 2230
rect 12560 1618 12570 2230
rect 12600 1546 12724 2390
rect 12856 2386 13542 2390
rect 12754 1618 12764 2230
rect 12818 1618 12828 2230
rect 12856 1546 12982 2386
rect 13012 1618 13022 2230
rect 13076 1618 13086 2230
rect 13294 1454 13300 1457
rect 6907 1408 13300 1454
rect 6820 632 6830 1244
rect 6884 632 6894 1244
rect 6924 560 7048 1408
rect 7078 630 7088 1242
rect 7142 630 7152 1242
rect 7182 560 7306 1408
rect 7336 632 7346 1244
rect 7400 632 7410 1244
rect 7440 472 7564 1316
rect 7594 632 7604 1244
rect 7658 632 7668 1244
rect 7698 472 7822 1316
rect 7852 632 7862 1244
rect 7916 632 7926 1244
rect 7956 472 8080 1316
rect 8110 632 8120 1244
rect 8174 632 8184 1244
rect 8214 472 8338 1316
rect 8368 632 8378 1244
rect 8432 632 8442 1244
rect 8472 560 8596 1408
rect 8732 1316 8856 1408
rect 8730 1270 8856 1316
rect 8626 632 8636 1244
rect 8690 632 8700 1244
rect 8730 560 8854 1270
rect 8884 632 8894 1244
rect 8948 632 8958 1244
rect 8988 560 9112 1408
rect 9142 632 9152 1244
rect 9206 632 9216 1244
rect 9246 560 9370 1408
rect 9400 632 9410 1244
rect 9464 632 9474 1244
rect 9504 472 9628 1316
rect 9658 632 9668 1244
rect 9722 632 9732 1244
rect 9762 472 9886 1316
rect 9916 632 9926 1246
rect 9978 632 9988 1246
rect 10020 472 10144 1316
rect 10174 632 10184 1244
rect 10238 632 10248 1244
rect 10278 472 10402 1316
rect 10432 632 10442 1244
rect 10496 632 10506 1244
rect 10536 560 10660 1408
rect 10690 632 10700 1244
rect 10754 632 10764 1244
rect 10794 560 10918 1408
rect 10948 632 10958 1244
rect 11012 632 11022 1244
rect 11052 560 11176 1408
rect 11206 632 11216 1244
rect 11270 632 11280 1244
rect 11310 560 11434 1408
rect 11464 632 11474 1244
rect 11528 632 11538 1244
rect 11568 472 11692 1316
rect 11722 632 11732 1244
rect 11786 632 11796 1244
rect 11826 472 11950 1316
rect 11980 632 11990 1244
rect 12044 632 12054 1244
rect 12084 472 12208 1316
rect 12238 632 12248 1244
rect 12302 632 12312 1244
rect 12342 472 12466 1316
rect 12496 632 12506 1244
rect 12560 632 12570 1244
rect 12600 560 12724 1408
rect 12754 632 12764 1244
rect 12818 632 12828 1244
rect 12858 560 12982 1408
rect 13294 1405 13300 1408
rect 13352 1405 13358 1457
rect 13012 632 13022 1244
rect 13076 632 13086 1244
rect 13474 472 13542 2386
rect 7416 404 13542 472
rect 6287 276 6357 282
rect 5518 166 5570 172
rect 5518 108 5570 114
rect 7895 166 7947 172
rect 7895 108 7947 114
rect 5316 104 5326 106
rect 5256 -108 5266 104
rect 5438 -10 5448 106
rect 5822 -2 5832 64
rect 6914 -2 6924 64
rect 7896 54 7946 108
rect 10965 103 11067 109
rect 7380 4 8462 54
rect 5370 -16 5434 -10
rect 5370 -108 5381 -16
rect 4918 -490 4994 -484
rect 5094 -670 5146 -664
rect 5094 -728 5146 -722
rect 3950 -2164 3992 -1230
rect 4736 -1300 4746 -1054
rect 4822 -1300 4832 -1054
rect 4756 -1519 4808 -1300
rect 4944 -1359 4950 -1282
rect 5027 -1359 5033 -1282
rect 4732 -1525 4809 -1519
rect 4732 -1608 4809 -1602
rect 4950 -1525 5027 -1359
rect 4950 -1608 5027 -1602
rect 3016 -2232 3026 -2178
rect 3080 -2232 3090 -2178
rect 930 -3290 948 -3204
rect 1042 -3290 1060 -3204
rect 1382 -3202 1512 -2350
rect 1382 -3288 1398 -3202
rect 1492 -3288 1512 -3202
rect 1382 -3290 1512 -3288
rect 1842 -3204 1972 -2350
rect 2114 -2850 2160 -2238
rect 1842 -3290 1856 -3204
rect 1950 -3290 1972 -3204
rect 2298 -3202 2428 -2350
rect 2298 -3288 2314 -3202
rect 2408 -3288 2428 -3202
rect 2298 -3290 2428 -3288
rect 2756 -3204 2886 -2352
rect 3030 -2842 3076 -2232
rect 3932 -2244 3942 -2164
rect 4022 -2244 4032 -2164
rect 3950 -2246 3992 -2244
rect 4366 -2536 4492 -2462
rect 4756 -2536 4808 -1608
rect 4366 -2614 4808 -2536
rect 4366 -2690 4688 -2614
rect 4798 -2690 4808 -2614
rect 5095 -2620 5145 -728
rect 5094 -2626 5146 -2620
rect 5094 -2684 5146 -2678
rect 4366 -2846 4808 -2690
rect 4366 -2920 4492 -2846
rect 5304 -2962 5381 -108
rect 5832 -1048 5882 -2
rect 5920 -1068 6052 -62
rect 5910 -1120 5920 -1068
rect 6052 -1120 6062 -1068
rect 6090 -1210 6140 -136
rect 6178 -1068 6310 -62
rect 6348 -1048 6398 -2
rect 6168 -1120 6178 -1068
rect 6310 -1120 6320 -1068
rect 6436 -1070 6568 -62
rect 6426 -1122 6436 -1070
rect 6568 -1122 6578 -1070
rect 6606 -1210 6656 -136
rect 6694 -1074 6826 -62
rect 6864 -1048 6914 -2
rect 7380 -1048 7430 4
rect 7468 -1064 7600 -62
rect 6684 -1130 6694 -1074
rect 6826 -1130 6836 -1074
rect 7458 -1120 7468 -1064
rect 7600 -1120 7610 -1064
rect 6090 -1264 6656 -1210
rect 7638 -1206 7688 -136
rect 7726 -1064 7858 -62
rect 7896 -1048 7946 4
rect 7984 -1064 8116 -62
rect 7716 -1120 7726 -1064
rect 7858 -1120 7868 -1064
rect 7974 -1120 7984 -1064
rect 8116 -1120 8126 -1064
rect 8154 -1206 8204 -136
rect 8242 -1064 8374 -62
rect 8412 -1048 8462 4
rect 8928 22 10965 82
rect 8928 -1048 8978 22
rect 9016 -1064 9148 -64
rect 8232 -1120 8242 -1064
rect 8374 -1120 8384 -1064
rect 9006 -1120 9016 -1064
rect 9148 -1120 9158 -1064
rect 7638 -1262 8206 -1206
rect 9186 -1214 9236 -136
rect 9274 -1064 9406 -64
rect 9444 -1048 9494 22
rect 9532 -1064 9664 -64
rect 9264 -1120 9274 -1064
rect 9406 -1120 9416 -1064
rect 9522 -1120 9532 -1064
rect 9664 -1120 9674 -1064
rect 9702 -1214 9752 -136
rect 9790 -1064 9922 -64
rect 9960 -1048 10010 22
rect 10048 -1064 10180 -64
rect 9780 -1120 9790 -1064
rect 9922 -1120 9932 -1064
rect 10038 -1120 10048 -1064
rect 10180 -1120 10190 -1064
rect 10218 -1214 10268 -136
rect 10306 -1064 10438 -64
rect 10476 -1048 10526 22
rect 11067 22 13106 82
rect 10965 -5 11067 1
rect 10564 -1064 10696 -64
rect 10296 -1120 10306 -1064
rect 10438 -1120 10448 -1064
rect 10554 -1120 10564 -1064
rect 10696 -1120 10706 -1064
rect 10734 -1214 10784 -136
rect 10822 -1064 10954 -64
rect 10992 -1050 11042 -5
rect 11080 -1064 11212 -64
rect 10812 -1120 10822 -1064
rect 10954 -1120 10964 -1064
rect 11070 -1120 11080 -1064
rect 11212 -1120 11222 -1064
rect 11250 -1214 11300 -136
rect 11338 -1064 11470 -64
rect 11508 -1048 11558 22
rect 11596 -1064 11728 -64
rect 11328 -1120 11338 -1064
rect 11470 -1120 11480 -1064
rect 11586 -1120 11596 -1064
rect 11728 -1120 11738 -1064
rect 11766 -1214 11816 -136
rect 11854 -1064 11986 -64
rect 12024 -1048 12074 22
rect 12112 -1064 12244 -64
rect 11844 -1120 11854 -1064
rect 11986 -1120 11996 -1064
rect 12102 -1120 12112 -1064
rect 12244 -1120 12254 -1064
rect 12282 -1214 12332 -136
rect 12370 -1064 12502 -64
rect 12540 -1048 12590 22
rect 12628 -1064 12760 -64
rect 12360 -1120 12370 -1064
rect 12502 -1120 12512 -1064
rect 12618 -1120 12628 -1064
rect 12760 -1120 12770 -1064
rect 12798 -1214 12848 -136
rect 12886 -1064 13018 -64
rect 13056 -1048 13106 22
rect 13526 -758 13598 -752
rect 13526 -836 13598 -830
rect 12876 -1120 12886 -1064
rect 13018 -1120 13028 -1064
rect 7638 -1264 7688 -1262
rect 6208 -1622 6260 -1616
rect 6208 -1680 6260 -1674
rect 5280 -3040 5384 -2962
rect 5280 -3146 5290 -3040
rect 5482 -3146 5492 -3040
rect 2756 -3290 2770 -3204
rect 2864 -3290 2886 -3204
rect 930 -3292 1060 -3290
rect 2756 -3292 2886 -3290
rect -3955 -3306 -3845 -3300
rect -4132 -3516 -4080 -3510
rect 5320 -3458 5372 -3146
rect 5320 -3516 5372 -3510
rect -4267 -3603 -4213 -3597
rect 6211 -3914 6257 -1680
rect 6319 -3108 6389 -1264
rect 6814 -1686 6824 -1614
rect 6890 -1686 6900 -1614
rect 7330 -1686 7340 -1614
rect 7406 -1686 7416 -1614
rect 7846 -1686 7856 -1614
rect 7922 -1686 7932 -1614
rect 6832 -2848 6882 -1686
rect 6920 -3064 7052 -1864
rect 7178 -3064 7310 -1864
rect 7348 -2848 7398 -1686
rect 7436 -3064 7568 -1864
rect 7694 -3064 7826 -1864
rect 7864 -2848 7914 -1686
rect 8154 -1734 8204 -1262
rect 9186 -1264 12848 -1214
rect 8878 -1686 8888 -1614
rect 8954 -1686 8964 -1614
rect 9910 -1686 9920 -1614
rect 9986 -1686 9996 -1614
rect 10942 -1686 10952 -1614
rect 11018 -1686 11028 -1614
rect 11746 -1618 11818 -1264
rect 13527 -1286 13598 -836
rect 13527 -1363 13598 -1357
rect 13660 -1386 13712 2770
rect 13788 2686 13843 2692
rect 13788 -1224 13843 2631
rect 14701 2474 14751 3432
rect 15618 3384 15670 3390
rect 13920 2468 13972 2474
rect 13920 2410 13972 2416
rect 14700 2468 14752 2474
rect 14700 2410 14752 2416
rect 13921 696 13971 2410
rect 15618 2294 15670 3332
rect 16577 2430 16627 3433
rect 16718 3432 16768 3433
rect 16576 2424 16628 2430
rect 16576 2366 16628 2372
rect 17272 2294 17320 4770
rect 19200 4766 19252 4772
rect 18106 4600 18186 4606
rect 18750 4522 18760 4574
rect 18884 4522 19018 4574
rect 19142 4522 19276 4574
rect 19400 4522 19534 4574
rect 19658 4522 19668 4574
rect 18106 3114 18186 4520
rect 18668 3517 18718 4494
rect 18760 3600 18884 4522
rect 18926 3680 18976 4522
rect 19018 3600 19142 4522
rect 19184 3517 19234 4494
rect 19276 3600 19400 4522
rect 19442 3680 19492 4522
rect 19534 3600 19658 4522
rect 19700 3517 19750 4494
rect 20308 3652 20432 4574
rect 20474 3652 20524 4494
rect 20566 3652 20690 4574
rect 20731 3652 20781 3655
rect 20824 3652 20948 4574
rect 20990 3652 21040 4494
rect 21082 3652 21206 4574
rect 20298 3600 20308 3652
rect 20432 3600 20566 3652
rect 20690 3600 20824 3652
rect 20948 3600 21082 3652
rect 21206 3600 21216 3652
rect 20731 3517 20781 3600
rect 18668 3467 20781 3517
rect 21853 3557 21932 3563
rect 21702 3344 21774 3350
rect 18106 3028 18186 3034
rect 18923 3277 18981 3283
rect 17690 2424 17742 2430
rect 17690 2366 17742 2372
rect 17911 2421 17977 2427
rect 14692 2242 15772 2294
rect 16754 2250 17320 2294
rect 14514 2090 14524 2142
rect 14652 2090 14662 2142
rect 14434 1490 14482 2064
rect 14524 1580 14652 2090
rect 14692 1654 14740 2242
rect 14772 2090 14782 2142
rect 14910 2090 14920 2142
rect 15030 2090 15040 2142
rect 15168 2090 15178 2142
rect 14782 1580 14910 2090
rect 14950 1490 14998 2066
rect 15040 1580 15168 2090
rect 15208 1654 15256 2242
rect 15288 2090 15298 2142
rect 15426 2090 15436 2142
rect 15546 2090 15556 2142
rect 15684 2090 15694 2142
rect 15298 1580 15426 2090
rect 15466 1490 15514 2066
rect 15556 1580 15684 2090
rect 15724 1654 15772 2242
rect 15804 2090 15814 2142
rect 15942 2090 15952 2142
rect 16578 2090 16588 2142
rect 16718 2090 16728 2142
rect 15814 1580 15942 2090
rect 15982 1490 16030 2066
rect 14432 1436 16030 1490
rect 16498 1496 16546 2066
rect 16588 1580 16718 2090
rect 16756 1654 16804 2250
rect 16836 2090 16846 2142
rect 16976 2090 16986 2142
rect 17092 2090 17102 2142
rect 17232 2090 17242 2142
rect 16846 1580 16976 2090
rect 17014 1496 17062 2066
rect 17102 1580 17232 2090
rect 17272 1654 17320 2250
rect 16498 1438 17062 1496
rect 13920 690 13972 696
rect 15140 692 15226 1436
rect 16728 1035 16802 1438
rect 17691 1018 17741 2366
rect 17911 2147 17977 2355
rect 18923 2266 18981 3219
rect 17911 2075 17977 2081
rect 18532 2144 19614 2266
rect 18532 2090 18624 2144
rect 18748 2104 19614 2144
rect 18748 2090 18758 2104
rect 18882 2090 19264 2104
rect 18532 1652 18582 2090
rect 18624 1580 18748 2090
rect 18790 1484 18840 2064
rect 18882 1580 19006 2090
rect 19048 1652 19098 2090
rect 19140 1580 19264 2090
rect 19398 2090 19614 2104
rect 19306 1484 19356 2064
rect 19398 1580 19522 2090
rect 19564 1652 19614 2090
rect 20172 1630 20296 2136
rect 20338 1630 20388 2064
rect 20430 1630 20554 2136
rect 20170 1628 20554 1630
rect 20688 1628 20812 2136
rect 20854 1628 20904 2064
rect 20946 1628 21070 2136
rect 20168 1570 21074 1628
rect 20338 1484 20388 1570
rect 20854 1484 20904 1570
rect 18790 1436 20904 1484
rect 19581 1035 19655 1041
rect 16728 955 16802 961
rect 17690 1012 17742 1018
rect 17690 954 17742 960
rect 15920 878 15992 884
rect 15920 692 15992 806
rect 19581 694 19655 961
rect 21580 878 21652 884
rect 13920 632 13972 638
rect 14432 690 17578 692
rect 14432 644 15166 690
rect 14432 -748 14482 644
rect 14524 -768 14648 536
rect 14514 -820 14524 -768
rect 14648 -820 14658 -768
rect 14690 -894 14740 464
rect 14782 -768 14906 536
rect 14948 -748 14998 644
rect 15218 644 17578 690
rect 15166 632 15218 638
rect 15040 -768 15164 536
rect 14772 -820 14782 -768
rect 14906 -820 14916 -768
rect 15030 -820 15040 -768
rect 15164 -820 15174 -768
rect 15206 -894 15256 464
rect 15298 -768 15422 536
rect 15464 -748 15514 644
rect 15920 624 16030 644
rect 15556 -768 15680 536
rect 15288 -820 15298 -768
rect 15422 -820 15432 -768
rect 15546 -820 15556 -768
rect 15680 -820 15690 -768
rect 15722 -894 15772 464
rect 15814 -768 15938 536
rect 15980 -748 16030 624
rect 16072 -768 16196 536
rect 15804 -820 15814 -768
rect 15938 -820 15948 -768
rect 16062 -820 16072 -768
rect 16196 -820 16206 -768
rect 16238 -894 16288 464
rect 16330 -768 16454 536
rect 16496 -748 16546 644
rect 16588 -768 16712 536
rect 16320 -820 16330 -768
rect 16454 -820 16464 -768
rect 16578 -820 16588 -768
rect 16712 -820 16722 -768
rect 16754 -894 16804 464
rect 16846 -768 16970 536
rect 17012 -748 17062 644
rect 17104 -768 17228 536
rect 16836 -820 16846 -768
rect 16970 -820 16980 -768
rect 17094 -820 17104 -768
rect 17228 -820 17238 -768
rect 17270 -894 17320 464
rect 17362 -768 17486 536
rect 17528 -748 17578 644
rect 18044 646 21190 694
rect 18044 -748 18094 646
rect 18136 -768 18260 536
rect 17352 -820 17362 -768
rect 17486 -820 17496 -768
rect 18126 -820 18136 -768
rect 18260 -820 18270 -768
rect 14690 -964 17320 -894
rect 18302 -908 18352 464
rect 18394 -768 18518 536
rect 18560 -748 18610 646
rect 18652 -768 18776 536
rect 18384 -820 18394 -768
rect 18518 -820 18528 -768
rect 18642 -820 18652 -768
rect 18776 -820 18786 -768
rect 18818 -908 18868 464
rect 18910 -768 19034 536
rect 19076 -748 19126 646
rect 19168 -768 19292 536
rect 18900 -820 18910 -768
rect 19034 -820 19044 -768
rect 19158 -820 19168 -768
rect 19292 -820 19302 -768
rect 19334 -908 19384 464
rect 19426 -768 19550 536
rect 19592 -748 19642 646
rect 19684 -768 19808 536
rect 19416 -820 19426 -768
rect 19550 -820 19560 -768
rect 19674 -820 19684 -768
rect 19808 -820 19818 -768
rect 19850 -908 19900 464
rect 19942 -768 20066 536
rect 20108 -750 20158 646
rect 20200 -768 20324 536
rect 19932 -820 19942 -768
rect 20066 -820 20076 -768
rect 20190 -820 20200 -768
rect 20324 -820 20334 -768
rect 20366 -908 20416 464
rect 20458 -768 20582 536
rect 20624 -748 20674 646
rect 20716 -768 20840 536
rect 20448 -820 20458 -768
rect 20582 -820 20592 -768
rect 20706 -820 20716 -768
rect 20840 -820 20850 -768
rect 20882 -908 20932 464
rect 20974 -768 21098 536
rect 21140 -748 21190 646
rect 20964 -820 20974 -768
rect 21098 -820 21108 -768
rect 18302 -964 20932 -908
rect 13982 -1218 14034 -1212
rect 14678 -1270 14688 -1218
rect 14742 -1270 14752 -1218
rect 13982 -1276 14034 -1270
rect 13788 -1285 13843 -1279
rect 13660 -1444 13712 -1438
rect 11670 -1686 11680 -1618
rect 11882 -1686 11892 -1618
rect 11974 -1686 11984 -1614
rect 12050 -1686 12060 -1614
rect 12490 -1686 12500 -1614
rect 12566 -1686 12576 -1614
rect 13006 -1686 13016 -1614
rect 13082 -1686 13092 -1614
rect 8138 -1800 8148 -1734
rect 8406 -1738 8416 -1734
rect 8432 -1790 8442 -1738
rect 8406 -1800 8430 -1790
rect 7952 -3064 8084 -1864
rect 8210 -3064 8342 -1864
rect 8380 -2848 8430 -1800
rect 8468 -3064 8600 -1864
rect 8726 -3064 8858 -1864
rect 8896 -2848 8946 -1686
rect 8984 -3064 9116 -1864
rect 9242 -3064 9374 -1864
rect 6318 -3188 6390 -3108
rect 6910 -3124 6920 -3064
rect 9364 -3124 9374 -3064
rect 9242 -3134 9374 -3124
rect 9412 -3188 9462 -1936
rect 9500 -3064 9632 -1864
rect 9758 -3064 9890 -1864
rect 9928 -2850 9978 -1686
rect 10016 -3064 10148 -1864
rect 10274 -3054 10406 -1864
rect 10274 -3064 10408 -3054
rect 9500 -3124 9510 -3064
rect 10396 -3124 10408 -3064
rect 9500 -3134 9632 -3124
rect 10274 -3136 10408 -3124
rect 10444 -3188 10494 -1936
rect 10532 -3064 10664 -1864
rect 10790 -3064 10922 -1864
rect 10960 -2850 11010 -1686
rect 11464 -1786 11474 -1734
rect 11528 -1786 11538 -1734
rect 11048 -3064 11180 -1864
rect 11306 -3064 11438 -1864
rect 11476 -2848 11526 -1786
rect 11564 -3064 11696 -1864
rect 11822 -3064 11954 -1864
rect 11992 -2848 12042 -1686
rect 12080 -3064 12212 -1864
rect 12338 -3064 12470 -1864
rect 12508 -2848 12558 -1686
rect 12596 -3064 12728 -1864
rect 12854 -3064 12986 -1864
rect 13024 -2848 13074 -1686
rect 10532 -3124 10546 -3064
rect 12986 -3124 12996 -3064
rect 10532 -3134 10664 -3124
rect 6316 -3250 6326 -3188
rect 6388 -3250 6398 -3188
rect 9400 -3240 9410 -3188
rect 9464 -3240 9474 -3188
rect 10432 -3240 10442 -3188
rect 10496 -3240 10506 -3188
rect 13665 -3704 13711 -1444
rect 13662 -3710 13714 -3704
rect 13662 -3768 13714 -3762
rect 13987 -3818 14029 -1276
rect 14524 -2920 14648 -1564
rect 14690 -2848 14740 -1270
rect 15956 -1378 16056 -964
rect 19534 -1208 19676 -964
rect 16226 -1270 16236 -1218
rect 16290 -1270 16300 -1218
rect 16742 -1270 16752 -1218
rect 16806 -1270 16816 -1218
rect 18290 -1270 18300 -1218
rect 18354 -1270 18364 -1218
rect 18806 -1270 18816 -1218
rect 18870 -1270 18880 -1218
rect 15194 -1436 15204 -1384
rect 15258 -1436 15268 -1384
rect 15710 -1436 15720 -1384
rect 15774 -1436 15784 -1384
rect 14682 -2920 14737 -2919
rect 14782 -2920 14906 -1564
rect 15040 -2920 15164 -1564
rect 15206 -2848 15256 -1436
rect 15298 -2920 15422 -1564
rect 15556 -2920 15680 -1564
rect 15722 -2848 15772 -1436
rect 15914 -1450 15924 -1378
rect 16076 -1450 16086 -1378
rect 15814 -2920 15938 -1564
rect 16072 -2920 16196 -1564
rect 16238 -2848 16288 -1270
rect 16330 -2920 16454 -1564
rect 16588 -2920 16712 -1564
rect 16754 -2848 16804 -1270
rect 17258 -1436 17268 -1384
rect 17322 -1436 17332 -1384
rect 17774 -1436 17784 -1384
rect 17838 -1436 17848 -1384
rect 16846 -2920 16970 -1564
rect 17104 -2920 17228 -1564
rect 17270 -2848 17320 -1436
rect 17362 -2920 17486 -1564
rect 17620 -2920 17744 -1564
rect 17786 -2848 17836 -1436
rect 17878 -2920 18002 -1564
rect 18136 -2920 18260 -1564
rect 18302 -2848 18352 -1270
rect 18394 -2920 18518 -1564
rect 18652 -2920 18776 -1564
rect 18818 -2848 18868 -1270
rect 19508 -1280 19518 -1208
rect 19698 -1280 19708 -1208
rect 20354 -1270 20364 -1218
rect 20418 -1270 20428 -1218
rect 19322 -1436 19332 -1384
rect 19386 -1436 19396 -1384
rect 19836 -1436 19846 -1384
rect 19900 -1436 19910 -1384
rect 18910 -2920 19034 -1564
rect 19168 -2920 19292 -1564
rect 19334 -2848 19384 -1436
rect 19426 -2920 19550 -1564
rect 19684 -2920 19808 -1564
rect 19848 -2848 19898 -1436
rect 19942 -2920 20066 -1564
rect 20200 -2920 20324 -1564
rect 20366 -2848 20416 -1270
rect 20458 -2920 20582 -1564
rect 21580 -2910 21652 806
rect 21702 -814 21774 3272
rect 21853 -677 21932 3478
rect 22030 3344 22102 11846
rect 22200 3557 22279 12146
rect 22720 12225 23094 12231
rect 22799 12146 23094 12225
rect 22720 12140 23094 12146
rect 22584 12066 22656 12072
rect 22727 12066 23094 12140
rect 22578 11994 23094 12066
rect 22584 11864 22656 11994
rect 22727 11943 23094 11994
rect 22970 11856 23094 11943
rect 22584 11786 22656 11792
rect 22708 11367 22771 11373
rect 22402 9548 22454 9554
rect 22402 9490 22454 9496
rect 22403 8280 22453 9490
rect 22555 9428 22621 9435
rect 22555 9376 22562 9428
rect 22614 9376 22621 9428
rect 22402 8274 22454 8280
rect 22402 8216 22454 8222
rect 22200 3472 22279 3478
rect 22030 3266 22102 3272
rect 22028 3114 22108 3120
rect 22028 -528 22108 3034
rect 22555 2421 22621 9376
rect 22708 8169 22771 11304
rect 23339 11133 23400 14039
rect 23339 11066 23400 11072
rect 23461 13899 23519 13905
rect 23461 11004 23519 13841
rect 23589 13755 23655 13761
rect 23589 11749 23655 13689
rect 24136 11748 24260 12670
rect 24126 11696 24136 11748
rect 24260 11696 24270 11748
rect 23589 11677 23655 11683
rect 24304 11631 24350 12590
rect 24394 11748 24518 12670
rect 24652 11748 24776 12670
rect 24384 11696 24394 11748
rect 24518 11696 24528 11748
rect 24642 11696 24652 11748
rect 24776 11696 24786 11748
rect 24304 11598 24351 11631
rect 24305 11322 24351 11598
rect 24820 11322 24866 12590
rect 25336 11631 25382 12590
rect 25426 11748 25550 12670
rect 25684 11748 25808 12670
rect 25416 11696 25426 11748
rect 25550 11696 25560 11748
rect 25674 11696 25684 11748
rect 25808 11696 25818 11748
rect 25335 11598 25382 11631
rect 25335 11456 25381 11598
rect 25852 11456 25898 12590
rect 25942 11748 26066 12670
rect 26200 11748 26324 12670
rect 25932 11696 25942 11748
rect 26066 11696 26076 11748
rect 26190 11696 26200 11748
rect 26324 11696 26334 11748
rect 26368 11649 26414 12590
rect 26458 11748 26582 12670
rect 26716 11748 26840 12670
rect 26448 11696 26458 11748
rect 26582 11696 26592 11748
rect 26706 11696 26716 11748
rect 26840 11696 26850 11748
rect 26367 11572 26414 11649
rect 26884 11653 26930 12590
rect 26974 11748 27098 12670
rect 27232 11748 27356 12670
rect 26964 11696 26974 11748
rect 27098 11696 27108 11748
rect 27222 11696 27232 11748
rect 27356 11696 27366 11748
rect 26884 11602 26931 11653
rect 26882 11572 26931 11602
rect 26364 11566 26416 11572
rect 26364 11508 26416 11514
rect 26882 11566 26934 11572
rect 27400 11566 27446 12590
rect 27490 11748 27614 12670
rect 27748 11748 27872 12670
rect 27914 11748 27964 12590
rect 28006 11748 28130 12670
rect 28264 11748 28388 12670
rect 28430 11748 28480 12590
rect 28522 11748 28646 12670
rect 28780 11748 28904 12670
rect 28946 11748 28996 12590
rect 29038 11748 29162 12670
rect 29296 11748 29420 12670
rect 27480 11696 27490 11748
rect 27614 11696 27624 11748
rect 27738 11696 27748 11748
rect 28130 11696 28140 11748
rect 28254 11696 28264 11748
rect 28646 11696 28656 11748
rect 28770 11696 28780 11748
rect 29162 11696 29172 11748
rect 29286 11696 29296 11748
rect 29420 11696 29430 11748
rect 27914 11644 27964 11696
rect 28429 11658 28480 11696
rect 28946 11670 28996 11696
rect 28429 11593 28479 11658
rect 29462 11609 29512 12590
rect 29554 11748 29678 12670
rect 29812 11748 29936 12670
rect 29544 11696 29554 11748
rect 29678 11696 29688 11748
rect 29802 11696 29812 11748
rect 29936 11696 29946 11748
rect 27650 11568 27702 11574
rect 27391 11514 27397 11566
rect 27449 11514 27455 11566
rect 26882 11508 26934 11514
rect 27650 11510 27702 11516
rect 25332 11450 25384 11456
rect 25332 11392 25384 11398
rect 25849 11450 25901 11456
rect 25849 11392 25901 11398
rect 24302 11316 24354 11322
rect 24302 11258 24354 11264
rect 24451 11316 24503 11322
rect 24451 11258 24503 11264
rect 24817 11316 24869 11322
rect 24817 11258 24869 11264
rect 23428 10924 23438 11004
rect 23542 10924 23552 11004
rect 24452 10865 24502 11258
rect 27651 10871 27701 11510
rect 28430 11216 28478 11593
rect 29462 11572 29513 11609
rect 29462 11566 29516 11572
rect 29462 11564 29464 11566
rect 29464 11506 29516 11512
rect 29978 11570 30028 12590
rect 30070 11748 30194 12670
rect 30328 11748 30452 12670
rect 30060 11696 30070 11748
rect 30194 11696 30204 11748
rect 30318 11696 30328 11748
rect 30452 11696 30462 11748
rect 30494 11570 30544 12590
rect 30586 11748 30710 12670
rect 30844 11748 30968 12668
rect 30576 11696 30586 11748
rect 30710 11696 30720 11748
rect 30834 11696 30844 11748
rect 30968 11696 30978 11748
rect 30844 11694 30968 11696
rect 29978 11564 30030 11570
rect 29978 11506 30030 11512
rect 30494 11564 30546 11570
rect 31010 11564 31060 12590
rect 31102 11748 31226 12668
rect 31360 11748 31484 12668
rect 31092 11696 31102 11748
rect 31226 11696 31236 11748
rect 31350 11696 31360 11748
rect 31484 11696 31494 11748
rect 31102 11694 31226 11696
rect 31360 11694 31484 11696
rect 31526 11564 31576 12590
rect 32044 11625 32090 12590
rect 32134 11748 32258 12670
rect 32392 11748 32516 12670
rect 32124 11696 32134 11748
rect 32258 11696 32268 11748
rect 32382 11696 32392 11748
rect 32516 11696 32526 11748
rect 32560 11653 32606 12590
rect 32650 11748 32774 12670
rect 32640 11696 32650 11748
rect 32774 11696 32784 11748
rect 32044 11598 32091 11625
rect 30494 11506 30546 11512
rect 31011 11456 31057 11564
rect 29611 11450 29663 11456
rect 29611 11392 29663 11398
rect 31008 11450 31060 11456
rect 31527 11454 31573 11564
rect 28428 11210 28480 11216
rect 28428 11152 28480 11158
rect 29614 11139 29660 11392
rect 31008 11390 31060 11396
rect 31524 11448 31576 11454
rect 31524 11390 31576 11396
rect 32045 11322 32091 11598
rect 32559 11598 32606 11653
rect 32559 11322 32605 11598
rect 32042 11316 32094 11322
rect 32042 11258 32094 11264
rect 32556 11316 32608 11322
rect 32556 11258 32608 11264
rect 31676 11210 31728 11216
rect 31676 11152 31728 11158
rect 29611 11080 29672 11139
rect 29588 11067 29686 11080
rect 29588 11006 29605 11067
rect 29666 11006 29686 11067
rect 29588 10990 29686 11006
rect 29612 10875 29662 10990
rect 23420 10815 24503 10865
rect 25484 10862 28113 10871
rect 25484 10821 28114 10862
rect 23162 9703 23212 10670
rect 23254 9828 23378 10750
rect 23420 9858 23470 10815
rect 23512 9828 23636 10750
rect 23244 9776 23254 9828
rect 23378 9776 23388 9828
rect 23502 9776 23512 9828
rect 23636 9776 23646 9828
rect 23678 9703 23728 10670
rect 23770 9828 23894 10750
rect 23936 9858 23986 10815
rect 24028 9828 24152 10750
rect 23760 9776 23770 9828
rect 23894 9776 23904 9828
rect 24018 9776 24028 9828
rect 24152 9776 24162 9828
rect 24194 9703 24244 10670
rect 24286 9828 24410 10750
rect 24452 9858 24502 10815
rect 24544 9828 24668 10750
rect 24276 9776 24286 9828
rect 24410 9776 24420 9828
rect 24534 9776 24544 9828
rect 24668 9776 24678 9828
rect 24710 9703 24760 10670
rect 25226 9711 25276 10670
rect 25318 9828 25442 10750
rect 25484 9858 25534 10821
rect 25576 9828 25700 10750
rect 25308 9776 25318 9828
rect 25442 9776 25452 9828
rect 25566 9776 25576 9828
rect 25700 9776 25710 9828
rect 25742 9711 25792 10670
rect 25834 9828 25958 10750
rect 26000 9858 26050 10821
rect 26092 9828 26216 10750
rect 25824 9776 25834 9828
rect 25958 9776 25968 9828
rect 26082 9776 26092 9828
rect 26216 9776 26226 9828
rect 26258 9711 26308 10670
rect 26350 9828 26474 10750
rect 26516 9858 26566 10821
rect 26608 9828 26732 10750
rect 26340 9776 26350 9828
rect 26474 9776 26484 9828
rect 26598 9776 26608 9828
rect 26732 9776 26742 9828
rect 26774 9711 26824 10670
rect 26866 9828 26990 10750
rect 27032 9858 27082 10821
rect 27124 9828 27248 10750
rect 26856 9776 26866 9828
rect 26990 9776 27000 9828
rect 27114 9776 27124 9828
rect 27248 9776 27258 9828
rect 27290 9711 27340 10670
rect 27382 9828 27506 10750
rect 27548 9858 27598 10821
rect 27640 9828 27764 10750
rect 27372 9776 27382 9828
rect 27506 9776 27516 9828
rect 27630 9776 27640 9828
rect 27764 9776 27774 9828
rect 27806 9711 27856 10670
rect 27898 9828 28022 10750
rect 28064 9858 28114 10821
rect 29096 10825 30179 10875
rect 31678 10873 31726 11152
rect 31860 10873 32244 10874
rect 28156 9828 28280 10750
rect 27888 9776 27898 9828
rect 28022 9776 28032 9828
rect 28146 9776 28156 9828
rect 28280 9776 28290 9828
rect 28322 9711 28372 10670
rect 28838 9711 28888 10670
rect 28930 9828 29054 10750
rect 29096 9858 29146 10825
rect 29188 9828 29312 10750
rect 28920 9776 28930 9828
rect 29054 9776 29064 9828
rect 29178 9776 29188 9828
rect 29312 9776 29322 9828
rect 29354 9711 29404 10670
rect 29446 9828 29570 10750
rect 29612 9858 29662 10825
rect 29704 9828 29828 10750
rect 29436 9776 29446 9828
rect 29570 9776 29580 9828
rect 29694 9776 29704 9828
rect 29828 9776 29838 9828
rect 29870 9711 29920 10670
rect 29962 9828 30086 10750
rect 30128 9858 30178 10825
rect 31160 10823 32244 10873
rect 30220 9828 30344 10750
rect 29952 9776 29962 9828
rect 30086 9776 30096 9828
rect 30210 9776 30220 9828
rect 30344 9776 30354 9828
rect 30386 9711 30436 10670
rect 23162 9653 24761 9703
rect 25226 9661 28373 9711
rect 28838 9666 30436 9711
rect 30902 9713 30952 10670
rect 30994 9828 31118 10750
rect 31160 9858 31210 10823
rect 31252 9828 31376 10750
rect 31418 9828 31468 10670
rect 31510 9828 31634 10750
rect 31676 9858 31726 10823
rect 31860 10822 32244 10823
rect 31768 9828 31892 10750
rect 31934 9828 31984 10670
rect 32026 9828 32150 10750
rect 32192 9858 32242 10822
rect 32284 9828 32408 10750
rect 30984 9776 30994 9828
rect 32410 9776 32420 9828
rect 31418 9713 31468 9776
rect 31934 9716 31984 9776
rect 31920 9713 31996 9716
rect 32450 9713 32500 10670
rect 30902 9666 32500 9713
rect 28838 9661 30435 9666
rect 30902 9663 32499 9666
rect 23377 8422 23427 9653
rect 26481 9554 26531 9661
rect 26480 9548 26532 9554
rect 26480 9490 26532 9496
rect 29625 9434 29675 9661
rect 31920 9590 31996 9663
rect 31920 9508 31996 9514
rect 33326 9590 33402 9596
rect 29624 9428 29676 9434
rect 29624 9370 29676 9376
rect 23636 8712 23642 8784
rect 23714 8712 23720 8784
rect 24242 8722 24252 8774
rect 24376 8722 24386 8774
rect 24500 8722 24510 8774
rect 24634 8722 24644 8774
rect 24758 8722 24768 8774
rect 24892 8722 24902 8774
rect 25016 8722 25026 8774
rect 25150 8722 25160 8774
rect 25274 8722 25284 8774
rect 25408 8722 25418 8774
rect 25532 8722 25542 8774
rect 25666 8722 25676 8774
rect 25790 8722 25800 8774
rect 25924 8722 25934 8774
rect 26048 8722 26058 8774
rect 26182 8722 26192 8774
rect 26306 8722 26316 8774
rect 26440 8722 26450 8774
rect 26564 8722 26574 8774
rect 26698 8722 26708 8774
rect 26822 8722 26832 8774
rect 26956 8722 26966 8774
rect 27080 8722 27090 8774
rect 27214 8722 27224 8774
rect 27338 8722 27348 8774
rect 27472 8722 27482 8774
rect 27596 8722 27606 8774
rect 27730 8722 27740 8774
rect 27854 8722 27864 8774
rect 27988 8722 27998 8774
rect 28112 8722 28122 8774
rect 28246 8722 28256 8774
rect 28370 8722 28380 8774
rect 28504 8722 28514 8774
rect 28628 8722 28638 8774
rect 28762 8722 28772 8774
rect 28886 8722 28896 8774
rect 29020 8722 29030 8774
rect 29144 8722 29154 8774
rect 29278 8722 29288 8774
rect 29402 8722 29412 8774
rect 29536 8722 29546 8774
rect 29660 8722 29670 8774
rect 29794 8722 29804 8774
rect 29918 8722 29928 8774
rect 30052 8722 30062 8774
rect 30176 8722 30186 8774
rect 30310 8722 30320 8774
rect 30434 8722 30444 8774
rect 30568 8722 30578 8774
rect 30692 8722 30702 8774
rect 30826 8722 30836 8774
rect 30950 8722 30960 8774
rect 31084 8722 31094 8774
rect 31208 8722 31218 8774
rect 31342 8722 31352 8774
rect 31466 8722 31476 8774
rect 31600 8722 31610 8774
rect 31724 8722 31734 8774
rect 31858 8722 31868 8774
rect 31982 8722 31992 8774
rect 32116 8722 32126 8774
rect 32240 8722 32250 8774
rect 32374 8722 32384 8774
rect 23376 8416 23428 8422
rect 23376 8358 23428 8364
rect 22707 8160 22777 8169
rect 22707 8097 22708 8160
rect 22771 8097 22777 8160
rect 22707 4991 22777 8097
rect 22707 4915 22777 4921
rect 23642 4824 23714 8712
rect 23642 4746 23714 4752
rect 24252 3600 24376 8722
rect 24418 3522 24468 8700
rect 24510 3600 24634 8722
rect 24768 3600 24892 8722
rect 24934 3522 24984 8700
rect 25026 3600 25150 8722
rect 25284 3600 25408 8722
rect 25450 3522 25500 8700
rect 25542 3600 25666 8722
rect 25800 3600 25924 8722
rect 25966 3522 26016 8700
rect 26058 3600 26182 8722
rect 26316 3600 26440 8722
rect 26482 3522 26532 8700
rect 26574 3600 26698 8722
rect 26742 8675 26788 8687
rect 26742 3699 26748 8675
rect 26782 3699 26788 8675
rect 26742 3687 26788 3699
rect 26832 3600 26956 8722
rect 26998 3522 27048 8700
rect 27090 3600 27214 8722
rect 27348 3600 27472 8722
rect 27514 3522 27564 8700
rect 27606 3600 27730 8722
rect 27864 3600 27988 8722
rect 28030 3522 28080 8700
rect 28122 3600 28246 8722
rect 28380 3600 28504 8722
rect 28546 3522 28596 8700
rect 28638 3600 28762 8722
rect 28806 8675 28852 8687
rect 28806 3699 28812 8675
rect 28846 3699 28852 8675
rect 28806 3687 28852 3699
rect 28896 3600 29020 8722
rect 29062 3522 29112 8700
rect 29154 3600 29278 8722
rect 29412 3600 29536 8722
rect 29578 3522 29628 8700
rect 29670 3600 29794 8722
rect 29928 3600 30052 8722
rect 30094 3522 30144 8700
rect 30186 3600 30310 8722
rect 30444 3600 30568 8722
rect 30610 3522 30660 8700
rect 30702 3600 30826 8722
rect 30870 8675 30916 8687
rect 30870 3699 30876 8675
rect 30910 3699 30916 8675
rect 30870 3687 30916 3699
rect 30960 3600 31084 8722
rect 31126 3522 31176 8700
rect 31218 3600 31342 8722
rect 31476 3600 31600 8722
rect 31642 3522 31692 8700
rect 31734 3600 31858 8722
rect 31992 3600 32116 8722
rect 32158 3522 32208 8700
rect 32250 3600 32374 8722
rect 24400 3435 32229 3522
rect 22555 2349 22621 2355
rect 28302 2948 28718 3435
rect 28302 2666 28326 2948
rect 28650 2666 28718 2948
rect 28302 2114 28718 2666
rect 23162 2092 30952 2114
rect 23162 2032 30842 2092
rect 30902 2032 30952 2092
rect 23162 2008 30952 2032
rect 22419 1037 22505 1043
rect 22419 -340 22505 951
rect 22996 -350 23120 1886
rect 23162 -198 23212 2008
rect 23254 -350 23378 1886
rect 23512 -350 23636 1886
rect 23678 -198 23728 2008
rect 23770 -350 23894 1886
rect 24028 -350 24152 1886
rect 24194 -198 24244 2008
rect 24286 -350 24410 1886
rect 24544 -350 24668 1886
rect 24710 -198 24760 2008
rect 24802 -350 24926 1886
rect 25060 -350 25184 1886
rect 25226 -198 25276 2008
rect 25318 -350 25442 1886
rect 25576 -350 25700 1886
rect 25742 -198 25792 2008
rect 25834 -350 25958 1886
rect 26092 -350 26216 1886
rect 26258 -198 26308 2008
rect 26350 -350 26474 1886
rect 26608 -350 26732 1886
rect 26774 -198 26824 2008
rect 26866 -350 26990 1886
rect 27124 -350 27248 1886
rect 27290 -198 27340 2008
rect 27382 -350 27506 1886
rect 27640 -350 27764 1886
rect 27806 -198 27856 2008
rect 27898 -350 28022 1886
rect 28156 -350 28280 1886
rect 28322 -198 28372 2008
rect 28414 -350 28538 1886
rect 28672 -350 28796 1886
rect 28838 -198 28888 2008
rect 28930 -350 29054 1886
rect 29188 -350 29312 1886
rect 29354 -198 29404 2008
rect 29446 -350 29570 1886
rect 29704 -350 29828 1886
rect 29870 -198 29920 2008
rect 29962 -350 30086 1886
rect 30220 -350 30344 1886
rect 30386 -198 30436 2008
rect 30478 -350 30602 1886
rect 30736 -350 30860 1886
rect 30902 -198 30952 2008
rect 32006 2092 32066 2098
rect 30994 -350 31118 1886
rect 32006 1520 32066 2032
rect 32128 1520 32188 3435
rect 32714 2006 32810 2012
rect 32714 1904 32810 1910
rect 32734 1714 32790 1904
rect 32854 1750 32950 1756
rect 32734 1686 32798 1714
rect 32250 1624 32676 1654
rect 32250 1542 32310 1624
rect 32372 1542 32554 1570
rect 32616 1542 32676 1624
rect 32738 1520 32798 1686
rect 32854 1648 32950 1654
rect 32860 1520 32920 1648
rect 32006 -328 32066 -234
rect 32128 -282 32310 -232
rect 32372 -328 32432 -234
rect 22986 -416 22996 -350
rect 31120 -416 31130 -350
rect 32006 -358 32432 -328
rect 32494 -328 32554 -234
rect 32616 -282 32798 -232
rect 32860 -328 32920 -234
rect 32494 -358 32920 -328
rect 22419 -432 22505 -426
rect 22028 -614 22108 -608
rect 21853 -762 21932 -756
rect 21702 -824 21778 -814
rect 21774 -896 21778 -824
rect 21702 -902 21778 -896
rect 14514 -2972 14524 -2920
rect 20582 -2972 20592 -2920
rect 14682 -3542 14737 -2972
rect 21574 -2982 21580 -2910
rect 21652 -2982 21658 -2910
rect 14682 -3603 14737 -3597
rect 13982 -3824 14034 -3818
rect 13982 -3882 14034 -3876
rect 6208 -3920 6260 -3914
rect 6208 -3978 6260 -3972
rect 21705 -4029 21778 -902
rect 22532 -954 22582 -882
rect 23046 -954 23096 -882
rect 33326 -900 33402 9514
rect 23822 -910 23872 -900
rect 24338 -910 24388 -900
rect 24854 -910 24904 -900
rect 25370 -910 25420 -900
rect 25886 -910 25936 -900
rect 30014 -910 30064 -900
rect 30530 -910 30580 -900
rect 31046 -910 31096 -900
rect 31562 -910 31612 -900
rect 32078 -910 32128 -900
rect 22532 -996 23098 -954
rect 23812 -966 23822 -910
rect 25936 -966 25946 -910
rect 26908 -966 26918 -910
rect 29032 -966 29042 -910
rect 30004 -966 30014 -910
rect 32128 -966 32138 -910
rect 22532 -1550 22582 -996
rect 22618 -1058 22754 -996
rect 22876 -1058 23012 -996
rect 22614 -1110 22624 -1058
rect 22748 -1110 22758 -1058
rect 22872 -1110 22882 -1058
rect 23006 -1110 23016 -1058
rect 22618 -1622 22754 -1110
rect 22524 -1868 22534 -1796
rect 22600 -1868 22610 -1796
rect 21871 -1894 21923 -1888
rect 21871 -1952 21923 -1946
rect 21705 -4108 21778 -4102
rect 21876 -4209 21917 -1952
rect 22542 -2780 22592 -1868
rect 22788 -2287 22842 -1134
rect 22876 -1622 23012 -1110
rect 23046 -1550 23096 -996
rect 23646 -1110 23656 -1058
rect 23780 -1110 23790 -1058
rect 23564 -1690 23614 -1136
rect 23656 -1620 23780 -1110
rect 23822 -1548 23872 -966
rect 23904 -1110 23914 -1058
rect 24038 -1110 24048 -1058
rect 24162 -1110 24172 -1058
rect 24296 -1110 24306 -1058
rect 23912 -1620 24036 -1110
rect 24080 -1690 24130 -1136
rect 24172 -1620 24296 -1110
rect 24338 -1548 24388 -966
rect 24420 -1110 24430 -1058
rect 24554 -1110 24564 -1058
rect 24678 -1110 24688 -1058
rect 24812 -1110 24822 -1058
rect 24430 -1620 24554 -1110
rect 24596 -1690 24646 -1136
rect 24688 -1620 24812 -1110
rect 24854 -1550 24904 -966
rect 24936 -1110 24946 -1058
rect 25070 -1110 25080 -1058
rect 25194 -1110 25204 -1058
rect 25328 -1110 25338 -1058
rect 24946 -1620 25070 -1110
rect 25112 -1690 25162 -1136
rect 25204 -1620 25328 -1110
rect 25370 -1548 25420 -966
rect 25452 -1110 25462 -1058
rect 25586 -1110 25596 -1058
rect 25708 -1110 25718 -1058
rect 25842 -1110 25852 -1058
rect 25462 -1620 25586 -1110
rect 25628 -1690 25678 -1136
rect 25720 -1620 25844 -1110
rect 25886 -1548 25936 -966
rect 25968 -1110 25978 -1058
rect 26102 -1110 26112 -1058
rect 26742 -1110 26752 -1058
rect 26876 -1110 26886 -1058
rect 25978 -1620 26102 -1110
rect 26144 -1690 26194 -1136
rect 23564 -1732 26194 -1690
rect 26660 -1698 26710 -1136
rect 26752 -1620 26876 -1110
rect 26918 -1548 26968 -966
rect 26998 -1110 27008 -1058
rect 27132 -1110 27142 -1058
rect 27258 -1110 27268 -1058
rect 27392 -1110 27402 -1058
rect 27010 -1620 27134 -1110
rect 27176 -1698 27226 -1136
rect 27268 -1620 27392 -1110
rect 27432 -1548 27482 -966
rect 27516 -1110 27526 -1058
rect 27650 -1110 27660 -1058
rect 27774 -1110 27784 -1058
rect 27908 -1110 27918 -1058
rect 27526 -1620 27650 -1110
rect 27692 -1698 27742 -1136
rect 27784 -1620 27908 -1110
rect 27950 -1548 28000 -966
rect 28032 -1110 28042 -1058
rect 28166 -1110 28176 -1058
rect 28290 -1110 28300 -1058
rect 28424 -1110 28434 -1058
rect 28042 -1620 28166 -1110
rect 28208 -1698 28258 -1136
rect 28300 -1620 28424 -1110
rect 28466 -1548 28516 -966
rect 28548 -1110 28558 -1058
rect 28682 -1110 28692 -1058
rect 28806 -1110 28816 -1058
rect 28940 -1110 28950 -1058
rect 28558 -1620 28682 -1110
rect 28724 -1698 28774 -1136
rect 28816 -1620 28940 -1110
rect 28982 -1548 29032 -966
rect 29064 -1110 29074 -1058
rect 29198 -1110 29208 -1058
rect 29838 -1110 29848 -1058
rect 29972 -1110 29982 -1058
rect 29074 -1620 29198 -1110
rect 29240 -1698 29290 -1136
rect 23040 -1868 23050 -1796
rect 23116 -1868 23126 -1796
rect 22633 -2341 23021 -2287
rect 22634 -2946 22758 -2341
rect 22892 -2946 23016 -2341
rect 23058 -2780 23108 -1868
rect 24588 -1950 24598 -1878
rect 24664 -1950 24674 -1878
rect 23556 -2064 23566 -1992
rect 23632 -2064 23642 -1992
rect 24072 -2064 24082 -1992
rect 24148 -2064 24158 -1992
rect 22634 -2952 23016 -2946
rect 23150 -2952 23274 -2296
rect 23408 -2952 23532 -2296
rect 23574 -2782 23624 -2064
rect 23666 -2952 23790 -2296
rect 23924 -2952 24048 -2296
rect 24090 -2782 24140 -2064
rect 24606 -2782 24656 -1950
rect 24854 -2000 24904 -1732
rect 26660 -1744 29290 -1698
rect 29756 -1696 29806 -1134
rect 29848 -1620 29972 -1110
rect 30014 -1548 30064 -966
rect 30096 -1110 30106 -1058
rect 30230 -1110 30240 -1058
rect 30354 -1110 30364 -1058
rect 30488 -1110 30498 -1058
rect 30106 -1620 30230 -1110
rect 30272 -1696 30322 -1134
rect 30364 -1620 30488 -1110
rect 30530 -1548 30580 -966
rect 30612 -1110 30622 -1058
rect 30746 -1110 30756 -1058
rect 30870 -1110 30880 -1058
rect 31004 -1110 31014 -1058
rect 30622 -1620 30746 -1110
rect 30788 -1696 30838 -1134
rect 30880 -1620 31004 -1110
rect 31046 -1550 31096 -966
rect 31128 -1110 31138 -1058
rect 31262 -1110 31272 -1058
rect 31386 -1110 31396 -1058
rect 31520 -1110 31530 -1058
rect 31138 -1620 31262 -1110
rect 31304 -1696 31354 -1134
rect 31396 -1620 31520 -1110
rect 31562 -1548 31612 -966
rect 31644 -1110 31654 -1058
rect 31778 -1110 31788 -1058
rect 31902 -1110 31912 -1058
rect 32036 -1110 32046 -1058
rect 31654 -1620 31778 -1110
rect 31820 -1696 31870 -1134
rect 31912 -1620 32036 -1110
rect 32078 -1548 32128 -966
rect 33326 -982 33402 -976
rect 32160 -1110 32170 -1058
rect 32294 -1110 32304 -1058
rect 32170 -1620 32294 -1110
rect 32336 -1696 32386 -1134
rect 29756 -1742 32386 -1696
rect 25620 -1864 25630 -1792
rect 25696 -1864 25706 -1792
rect 25104 -1950 25114 -1878
rect 25180 -1950 25190 -1878
rect 24840 -2052 24850 -2000
rect 24908 -2052 24918 -2000
rect 24696 -2952 24820 -2296
rect 24956 -2952 25080 -2296
rect 25122 -2782 25172 -1950
rect 25216 -2952 25340 -2296
rect 25474 -2952 25598 -2296
rect 25640 -2780 25686 -1864
rect 26136 -1950 26146 -1878
rect 26212 -1950 26222 -1878
rect 27950 -1898 28000 -1744
rect 31046 -1786 31096 -1742
rect 28718 -1858 28728 -1796
rect 28792 -1858 28802 -1796
rect 31030 -1848 31040 -1786
rect 31104 -1848 31114 -1786
rect 31298 -1854 31308 -1792
rect 31368 -1854 31378 -1792
rect 31814 -1854 31824 -1792
rect 31884 -1854 31894 -1792
rect 25730 -2952 25854 -2296
rect 25988 -2952 26112 -2296
rect 26156 -2778 26202 -1950
rect 27932 -1954 27942 -1898
rect 28010 -1954 28020 -1898
rect 28200 -1964 28210 -1902
rect 28274 -1964 28284 -1902
rect 26652 -2064 26662 -1992
rect 26728 -2064 26738 -1992
rect 22624 -3006 22634 -2952
rect 22758 -2953 22892 -2952
rect 22758 -3006 22817 -2953
rect 22752 -3008 22817 -3006
rect 22875 -3006 22892 -2953
rect 23016 -3006 23026 -2952
rect 23140 -3006 23150 -2952
rect 23274 -3006 23284 -2952
rect 23398 -3006 23408 -2952
rect 23532 -3006 23542 -2952
rect 23656 -3006 23666 -2952
rect 23790 -3006 23800 -2952
rect 23914 -3006 23924 -2952
rect 24048 -3006 24058 -2952
rect 24686 -3006 24696 -2952
rect 24820 -3006 24830 -2952
rect 24946 -3006 24956 -2952
rect 25080 -3006 25090 -2952
rect 25206 -3006 25216 -2952
rect 25340 -3006 25350 -2952
rect 25464 -3006 25474 -2952
rect 25598 -3006 25608 -2952
rect 25720 -3006 25730 -2952
rect 25854 -3006 25864 -2952
rect 25978 -3006 25988 -2952
rect 26112 -3006 26122 -2952
rect 26244 -2954 26368 -2298
rect 26506 -2954 26630 -2298
rect 26672 -2780 26718 -2064
rect 27686 -2082 27696 -2020
rect 27760 -2082 27770 -2020
rect 27164 -2164 27174 -2094
rect 27250 -2164 27260 -2094
rect 26762 -2954 26886 -2298
rect 27022 -2954 27146 -2298
rect 27188 -2954 27232 -2164
rect 27280 -2954 27404 -2298
rect 27538 -2954 27662 -2298
rect 27704 -2780 27750 -2082
rect 27794 -2954 27918 -2298
rect 22875 -3008 22926 -3006
rect 26234 -3008 26244 -2954
rect 26368 -3008 26378 -2954
rect 26496 -3008 26506 -2954
rect 26630 -3008 26640 -2954
rect 26752 -3008 26762 -2954
rect 26886 -3008 26896 -2954
rect 27012 -3008 27022 -2954
rect 27404 -3008 27414 -2954
rect 27528 -3008 27538 -2954
rect 27662 -3008 27672 -2954
rect 27784 -3008 27794 -2954
rect 27918 -3008 27928 -2954
rect 28054 -2956 28178 -2300
rect 28220 -2780 28266 -1964
rect 28310 -2954 28434 -2298
rect 28568 -2954 28692 -2298
rect 28736 -2780 28782 -1858
rect 29234 -1962 29244 -1900
rect 29304 -1962 29314 -1900
rect 29750 -1960 29760 -1898
rect 29820 -1960 29830 -1898
rect 28826 -2954 28950 -2298
rect 29084 -2954 29208 -2298
rect 29250 -2780 29300 -1962
rect 29342 -2954 29466 -2298
rect 29600 -2954 29724 -2298
rect 29766 -2780 29816 -1960
rect 30264 -2080 30274 -2018
rect 30338 -2080 30348 -2018
rect 30782 -2080 30792 -2018
rect 30856 -2080 30866 -2018
rect 30282 -2780 30332 -2080
rect 30374 -2952 30498 -2296
rect 30632 -2952 30756 -2296
rect 30798 -2780 30848 -2080
rect 30890 -2952 31014 -2296
rect 31148 -2952 31272 -2296
rect 31314 -2780 31364 -1854
rect 31406 -2952 31530 -2296
rect 31664 -2952 31788 -2296
rect 31828 -2780 31878 -1854
rect 28044 -3010 28054 -2956
rect 28178 -3010 28188 -2956
rect 28300 -3008 28310 -2954
rect 28434 -3008 28444 -2954
rect 28558 -3008 28568 -2954
rect 28692 -3008 28702 -2954
rect 28816 -3008 28826 -2954
rect 28950 -3008 28960 -2954
rect 29074 -3008 29084 -2954
rect 29208 -3008 29218 -2954
rect 29332 -3008 29342 -2954
rect 29466 -3008 29476 -2954
rect 29590 -3008 29600 -2954
rect 29724 -3008 29734 -2954
rect 30364 -3006 30374 -2952
rect 30498 -3006 30508 -2952
rect 30622 -3006 30632 -2952
rect 30756 -3006 30766 -2952
rect 30880 -3006 30890 -2952
rect 31014 -3006 31024 -2952
rect 31138 -3006 31148 -2952
rect 31272 -3006 31282 -2952
rect 31396 -3006 31406 -2952
rect 31530 -3006 31540 -2952
rect 31654 -3006 31664 -2952
rect 31788 -3006 31798 -2952
rect 21870 -4215 21922 -4209
rect 21870 -4273 21922 -4267
rect -5137 -4411 -5079 -4399
rect 22817 -4341 22875 -3011
rect 22817 -4405 22875 -4399
rect -6456 -4728 33408 -4634
rect -6456 -5596 -4414 -4728
rect 33248 -5596 33408 -4728
rect -6456 -5756 33408 -5596
<< via1 >>
rect -4182 14039 -4121 14100
rect -5332 13702 -5248 13786
rect -5614 5022 -5550 5086
rect -8186 4185 -8122 4249
rect -8903 3284 -8841 3346
rect -6000 2710 -5948 2762
rect 23339 14039 23400 14100
rect -3947 13841 -3889 13899
rect -3771 13689 -3705 13755
rect -3561 13473 -3499 13535
rect 17467 13473 17529 13535
rect -3445 13341 -3387 13399
rect 17191 13341 17249 13399
rect -3334 13198 -3266 13266
rect 16971 13199 17037 13265
rect -3208 13074 -3148 13134
rect 2782 12928 2834 12980
rect 11554 12928 11606 12980
rect 11808 12942 11880 13014
rect -2916 12772 -2856 12832
rect 2186 12772 2246 12832
rect -3080 12560 -3008 12632
rect -3080 8902 -3008 8974
rect -2324 12570 -2200 12622
rect -2066 12570 -1942 12622
rect -1808 12570 -1684 12622
rect -1550 12570 -1426 12622
rect -1292 12570 -1168 12622
rect -1034 12570 -910 12622
rect -776 12570 -652 12622
rect -518 12570 -394 12622
rect -260 12570 -136 12622
rect -2 12570 122 12622
rect 256 12570 380 12622
rect 514 12570 638 12622
rect 772 12570 896 12622
rect 1030 12570 1154 12622
rect 1288 12570 1412 12622
rect 1546 12570 1670 12622
rect 2186 12582 2246 12642
rect 2596 12436 2676 12516
rect 2418 9880 2470 9932
rect 2256 9750 2308 9802
rect -2913 8755 -2859 8809
rect -986 8920 -930 8976
rect -3208 8646 -3148 8706
rect -3334 8538 -3266 8606
rect -3445 8435 -3387 8493
rect -3561 8317 -3499 8379
rect -3771 8065 -3705 8131
rect -1607 8065 -1541 8131
rect -3947 7851 -3889 7909
rect -1755 7851 -1697 7909
rect -4182 7633 -4121 7694
rect -1918 7633 -1857 7694
rect -3812 6244 -3748 6308
rect -1607 7009 -1541 7075
rect -1755 6837 -1697 6895
rect -1581 6837 -1523 6895
rect -1918 6034 -1857 6095
rect -1760 6034 -1700 6094
rect -3812 5022 -3748 5086
rect -3162 5900 -3076 5964
rect -2198 5892 -2140 5958
rect -2922 5778 -2374 5836
rect -3254 4838 -3022 4904
rect -2844 4664 -2768 4728
rect -2274 4846 -2042 4912
rect -2528 4664 -2452 4728
rect -1581 5809 -1523 5867
rect -1760 4600 -1700 4660
rect -4028 4188 -3964 4252
rect -4210 3282 -4138 3354
rect -4562 2996 -4490 3068
rect -5178 2824 -5126 2876
rect -5398 2710 -5346 2762
rect -4798 2710 -4746 2762
rect -5846 1405 -5794 1457
rect -5178 1405 -5126 1457
rect -5889 612 -5831 670
rect -5137 612 -5079 670
rect -5850 -180 -5798 -128
rect -5236 -180 -5184 -128
rect -5803 -960 -5717 -874
rect -5365 -960 -5279 -874
rect -5880 -1761 -5828 -1709
rect -5479 -1766 -5417 -1704
rect -5875 -2533 -5823 -2481
rect -5584 -2533 -5532 -2481
rect -5876 -3337 -5824 -3285
rect -5690 -3337 -5638 -3285
rect -5474 -3762 -5422 -3710
rect -5584 -3876 -5532 -3824
rect -5690 -3972 -5638 -3920
rect -5358 -4102 -5285 -4029
rect -5236 -4268 -5184 -4216
rect -4430 2824 -4378 2876
rect -3864 2798 -3812 2850
rect -4028 2416 -3964 2480
rect -4210 1880 -4138 1952
rect -4430 1538 -4378 1590
rect -3670 2710 -3618 2762
rect -3502 2614 -3450 2666
rect -2671 2614 -2619 2666
rect -2914 2418 -2862 2470
rect -2428 2418 -2376 2470
rect -2756 1890 -2704 1942
rect -2586 1890 -2534 1942
rect 322 8646 382 8706
rect -533 8435 -475 8493
rect -653 8317 -591 8379
rect -913 7009 -847 7075
rect -595 5809 -537 5867
rect -986 4882 -926 4942
rect -1636 3268 -1580 3324
rect -1234 3268 -1178 3324
rect -1698 2904 -1644 2958
rect -1500 2798 -1448 2850
rect 433 8537 503 8607
rect 791 8479 853 8541
rect 796 7007 857 7068
rect 793 5807 851 5865
rect 364 3458 428 3522
rect -334 3268 -278 3324
rect 94 3268 150 3324
rect -592 3110 -540 3162
rect 806 4612 862 4668
rect 1894 8902 1966 8974
rect 1441 7293 1535 7387
rect 1689 8755 1743 8809
rect 1056 3268 1112 3324
rect 495 2731 561 2797
rect 1525 3219 1583 3277
rect -995 2645 -937 2703
rect -1500 1894 -1448 1946
rect -3185 1659 -3127 1717
rect -4582 1396 -4530 1448
rect -3864 1396 -3812 1448
rect 1525 1659 1583 1717
rect 1894 1754 1966 1826
rect 2090 8356 2166 8432
rect -2524 1538 -2472 1590
rect -4621 602 -4563 660
rect -3185 602 -3127 660
rect -4672 -162 -4618 -108
rect -4267 -162 -4213 -108
rect -4634 -844 -4582 -792
rect -4685 -1687 -4623 -1625
rect -4416 -2023 -4351 -1958
rect -4691 -3300 -4581 -3190
rect -3955 -521 -3881 -447
rect -4132 -844 -4080 -792
rect -3241 -521 -3167 -447
rect 1348 -502 1510 -448
rect -3740 -668 -3636 -588
rect -3241 -876 -3167 -802
rect -2336 -866 -2092 -812
rect -1878 -866 -1634 -812
rect -504 -866 -260 -812
rect -46 -866 198 -812
rect 412 -866 656 -812
rect 870 -866 1114 -812
rect 1328 -866 1572 -812
rect 1786 -866 2030 -812
rect -3584 -1036 -3458 -960
rect -3738 -1208 -3644 -1132
rect -3235 -1687 -3173 -1625
rect -3284 -1916 -3204 -1834
rect -2014 -1026 -1956 -970
rect -2474 -1904 -2412 -1844
rect -1558 -1904 -1496 -1844
rect -3736 -2356 -3640 -2264
rect -3100 -2023 -3035 -1958
rect -3107 -2244 -3029 -2166
rect -182 -1026 -124 -970
rect -2474 -2234 -2412 -2172
rect -1558 -2232 -1496 -2170
rect -642 -2232 -580 -2170
rect 734 -1026 792 -970
rect 1650 -1026 1708 -970
rect 9516 12582 9576 12642
rect 3396 12446 3520 12498
rect 3654 12446 3778 12498
rect 3912 12446 4036 12498
rect 4170 12446 4294 12498
rect 4428 12446 4552 12498
rect 4686 12446 4810 12498
rect 4944 12446 5068 12498
rect 5202 12446 5326 12498
rect 5460 12446 5584 12498
rect 5718 12446 5842 12498
rect 5976 12446 6100 12498
rect 6234 12446 6358 12498
rect 6492 12446 6616 12498
rect 6750 12446 6874 12498
rect 7008 12446 7132 12498
rect 7266 12446 7390 12498
rect 7524 12446 7648 12498
rect 7782 12446 7906 12498
rect 8040 12446 8164 12498
rect 8298 12446 8422 12498
rect 3560 10255 3614 10309
rect 4076 10253 4130 10307
rect 4592 10255 4646 10309
rect 5108 10255 5162 10309
rect 3799 10147 3853 10201
rect 6656 10253 6710 10307
rect 6888 10258 6940 10310
rect 7172 10255 7226 10309
rect 5883 10147 5937 10201
rect 9748 12448 9800 12500
rect 7688 10255 7742 10309
rect 9914 12448 10112 12500
rect 10230 12448 10428 12500
rect 10546 12448 10744 12500
rect 10862 12448 10914 12500
rect 12694 12946 12766 13018
rect 11808 12438 11880 12510
rect 14159 12883 14211 12935
rect 12308 12118 12398 12156
rect 12308 12046 12412 12118
rect 12308 12010 12398 12046
rect 12152 11768 12260 11850
rect 14675 12882 14727 12934
rect 15707 12881 15759 12933
rect 16223 12881 16275 12933
rect 15191 12739 15243 12791
rect 17191 12871 17249 12929
rect 16971 12049 17037 12115
rect 12976 11766 13084 11848
rect 11554 11494 11606 11546
rect 11810 11486 11926 11556
rect 20151 12873 20221 12943
rect 18348 12729 18420 12801
rect 18190 12056 18314 12108
rect 18448 12056 18572 12108
rect 19222 12056 19346 12108
rect 19480 12056 19604 12108
rect 19738 12056 19862 12108
rect 19996 12056 20120 12108
rect 20254 12056 20378 12108
rect 20512 12056 20636 12108
rect 20770 12056 20894 12108
rect 21028 12056 21152 12108
rect 22200 12146 22279 12225
rect 17467 11477 17529 11539
rect 18352 11494 18404 11546
rect 11684 11328 11756 11400
rect 11550 11158 11622 11230
rect 8203 10255 8257 10309
rect 9770 9880 9822 9932
rect 9554 9750 9606 9802
rect 3384 9486 3508 9538
rect 2780 8356 2856 8432
rect 2636 7428 2688 7480
rect 3642 9486 3766 9538
rect 3900 9486 4024 9538
rect 4158 9486 4282 9538
rect 4932 9486 5056 9538
rect 3812 7428 3864 7480
rect 5190 9486 5314 9538
rect 5448 9486 5572 9538
rect 5706 9486 5830 9538
rect 5964 9486 6088 9538
rect 6222 9486 6346 9538
rect 6480 9486 6604 9538
rect 6738 9486 6862 9538
rect 6996 9486 7120 9538
rect 6602 7388 6718 7504
rect 7254 9486 7378 9538
rect 7512 9486 7636 9538
rect 7770 9486 7894 9538
rect 8028 9486 8152 9538
rect 8286 9486 8410 9538
rect 8544 9486 8668 9538
rect 8802 9486 8926 9538
rect 9554 8364 9606 8416
rect 9770 8222 9822 8274
rect 10213 7401 10275 7463
rect 10898 8512 10977 8591
rect 10280 7146 10344 7210
rect 10138 6902 10190 6954
rect 2618 5792 2698 5876
rect 3254 5394 3310 6616
rect 3512 5394 3568 6616
rect 3770 5394 3826 6616
rect 4028 5394 4084 6616
rect 4286 5394 4342 6616
rect 4544 5394 4600 6616
rect 4802 5394 4858 6616
rect 5060 5394 5116 6616
rect 5318 5394 5374 6616
rect 5576 5394 5632 6616
rect 5834 5394 5890 6616
rect 6092 5394 6148 6616
rect 6350 5394 6406 6616
rect 6608 5394 6664 6616
rect 6866 5394 6922 6616
rect 7124 5394 7180 6616
rect 7382 5394 7438 6616
rect 7640 5394 7696 6616
rect 7898 5394 7954 6616
rect 8156 5394 8212 6616
rect 8414 5394 8470 6616
rect 8672 5394 8728 6616
rect 8930 5394 8986 6616
rect 9188 5394 9244 6616
rect 9446 5394 9502 6616
rect 3254 3790 3310 5012
rect 3512 3790 3568 5012
rect 3770 3790 3826 5012
rect 4028 3790 4084 5012
rect 4286 3790 4342 5012
rect 4544 3790 4600 5012
rect 4802 3790 4858 5012
rect 5060 3790 5116 5012
rect 5318 3790 5374 5012
rect 5576 3790 5632 5012
rect 5834 3790 5890 5012
rect 6092 3790 6148 5012
rect 6350 3790 6406 5012
rect 6608 3790 6664 5012
rect 6866 3790 6922 5012
rect 7124 3790 7180 5012
rect 7382 3790 7438 5012
rect 7640 3790 7696 5012
rect 7898 3790 7954 5012
rect 8156 3790 8212 5012
rect 8414 3790 8470 5012
rect 8672 3790 8728 5012
rect 8930 3790 8986 5012
rect 9188 3790 9244 5012
rect 9446 3790 9502 5012
rect 6041 3346 6120 3425
rect 2834 3004 2886 3056
rect 4760 1894 4812 1946
rect 3450 1754 3522 1826
rect 2636 1526 2688 1578
rect 2416 1380 2472 1436
rect 2902 -348 2958 -296
rect 3072 -348 3274 -296
rect 3100 -466 3220 -414
rect 3388 -348 3590 -296
rect 3704 -348 3906 -296
rect 4020 -348 4076 -296
rect 5518 1526 5570 1578
rect 5378 1380 5434 1436
rect 4898 876 5010 1186
rect 4748 -358 4820 -286
rect 3882 -476 4004 -418
rect 2256 -722 2308 -670
rect 2244 -866 2488 -812
rect 2702 -866 2946 -812
rect 3160 -866 3404 -812
rect 3618 -866 3862 -812
rect 2090 -1036 2166 -960
rect -3738 -2910 -3642 -2818
rect -3282 -3120 -3202 -3038
rect -3955 -3300 -3845 -3190
rect -2264 -3290 -2170 -3204
rect -1804 -3290 -1710 -3204
rect -1340 -3288 -1246 -3202
rect 256 -2242 352 -2174
rect 1190 -2232 1252 -2170
rect 2566 -1026 2624 -970
rect -886 -3280 -792 -3194
rect -432 -3290 -338 -3204
rect 260 -3108 348 -2962
rect 30 -3290 124 -3204
rect 482 -3292 576 -3206
rect 2106 -2238 2168 -2176
rect 3482 -1026 3540 -970
rect 10915 6997 10969 7051
rect 10449 5176 10507 5234
rect 10280 4918 10344 4982
rect 10138 3482 10190 3534
rect 10449 3477 10507 3535
rect 11184 8010 11256 8082
rect 11034 6904 11086 6956
rect 11684 9476 11756 9548
rect 19953 11304 20016 11367
rect 12314 11168 12438 11220
rect 12572 11168 12696 11220
rect 12830 11168 12954 11220
rect 13088 11168 13212 11220
rect 13346 11168 13470 11220
rect 13604 11168 13728 11220
rect 13862 11168 13986 11220
rect 14120 11168 14244 11220
rect 14378 11168 14502 11220
rect 14636 11168 14760 11220
rect 14894 11168 15018 11220
rect 15152 11168 15276 11220
rect 13666 8512 13745 8591
rect 15410 11168 15534 11220
rect 15668 11168 15792 11220
rect 15926 11168 16050 11220
rect 16184 11168 16308 11220
rect 16442 11168 16566 11220
rect 16700 11168 16824 11220
rect 16958 11168 17082 11220
rect 17216 11168 17340 11220
rect 17474 11168 17598 11220
rect 17732 11168 17856 11220
rect 17990 11168 18114 11220
rect 18248 11168 18372 11220
rect 18506 11168 18630 11220
rect 18764 11168 18888 11220
rect 19022 11168 19146 11220
rect 19280 11168 19404 11220
rect 19538 11168 19662 11220
rect 19796 11168 19920 11220
rect 20054 11168 20178 11220
rect 20312 11168 20436 11220
rect 20570 11168 20694 11220
rect 20828 11168 20952 11220
rect 21086 11168 21210 11220
rect 21344 11168 21468 11220
rect 11550 8010 11622 8082
rect 18683 8097 18746 8160
rect 11814 7886 11938 7938
rect 11184 5216 11256 5288
rect 12072 7886 12196 7938
rect 12330 7886 12454 7938
rect 12588 7886 12712 7938
rect 12846 7886 12970 7938
rect 13104 7886 13228 7938
rect 13362 7886 13486 7938
rect 13620 7886 13744 7938
rect 13878 7886 14002 7938
rect 14136 7886 14260 7938
rect 14394 7886 14518 7938
rect 14652 7886 14776 7938
rect 14910 7886 15034 7938
rect 11034 5066 11086 5118
rect 10898 3346 10977 3425
rect 9928 2846 9980 2898
rect 6041 1392 6120 1471
rect 6287 2483 6357 2553
rect 13144 5065 13199 5120
rect 12759 4921 12829 4991
rect 12560 4764 12612 4816
rect 12415 4519 12481 4585
rect 12560 3110 12612 3162
rect 12415 2731 12481 2797
rect 11195 2645 11253 2703
rect 12994 3482 13046 3534
rect 12994 2770 13046 2822
rect 14288 5216 14360 5288
rect 15168 7886 15292 7938
rect 15426 7886 15550 7938
rect 15684 7886 15808 7938
rect 15942 7886 16066 7938
rect 16200 7886 16324 7938
rect 16974 7886 17098 7938
rect 17232 7886 17356 7938
rect 17490 7886 17614 7938
rect 17748 7886 17872 7938
rect 18006 7886 18130 7938
rect 18264 7886 18388 7938
rect 18522 7886 18646 7938
rect 18780 7886 18904 7938
rect 19038 7886 19162 7938
rect 19296 7886 19420 7938
rect 19554 7886 19678 7938
rect 19812 7886 19936 7938
rect 20070 7886 20194 7938
rect 20328 7886 20452 7938
rect 20586 7886 20710 7938
rect 20844 7886 20968 7938
rect 21102 7886 21226 7938
rect 21360 7886 21484 7938
rect 16192 4772 16244 4824
rect 17270 4776 17322 4828
rect 19200 4772 19252 4824
rect 13972 4526 14096 4578
rect 14230 4526 14354 4578
rect 14488 4526 14612 4578
rect 14746 4526 14870 4578
rect 15004 4526 15128 4578
rect 15262 4526 15386 4578
rect 16036 4526 16160 4578
rect 16294 4526 16418 4578
rect 16552 4526 16676 4578
rect 13316 3332 13368 3384
rect 13144 2631 13199 2686
rect 13660 2770 13712 2822
rect 12759 2494 12829 2564
rect 6830 1618 6884 2230
rect 7088 1618 7142 2230
rect 7346 1618 7400 2230
rect 7604 1618 7658 2230
rect 7862 1618 7916 2230
rect 8120 1618 8174 2230
rect 8378 1618 8432 2230
rect 8636 1618 8690 2230
rect 8894 1618 8948 2230
rect 9152 1618 9206 2230
rect 9410 1618 9464 2230
rect 9668 1618 9722 2230
rect 9926 1618 9980 2230
rect 10184 1618 10238 2230
rect 10442 1618 10496 2230
rect 10700 1618 10754 2230
rect 10958 1618 11012 2230
rect 11216 1618 11270 2230
rect 11474 1618 11528 2230
rect 11732 1618 11786 2230
rect 11990 1618 12044 2230
rect 12248 1618 12302 2230
rect 12506 1618 12560 2230
rect 12764 1618 12818 2230
rect 13022 1618 13076 2230
rect 6830 632 6884 1244
rect 7088 630 7142 1242
rect 7346 632 7400 1244
rect 7604 632 7658 1244
rect 7862 632 7916 1244
rect 8120 632 8174 1244
rect 8378 632 8432 1244
rect 8636 632 8690 1244
rect 8894 632 8948 1244
rect 9152 632 9206 1244
rect 9410 632 9464 1244
rect 9668 632 9722 1244
rect 9926 632 9978 1246
rect 10184 632 10238 1244
rect 10442 632 10496 1244
rect 10700 632 10754 1244
rect 10958 632 11012 1244
rect 11216 632 11270 1244
rect 11474 632 11528 1244
rect 11732 632 11786 1244
rect 11990 632 12044 1244
rect 12248 632 12302 1244
rect 12506 632 12560 1244
rect 12764 632 12818 1244
rect 13300 1405 13352 1457
rect 13022 632 13076 1244
rect 6287 282 6357 352
rect 5518 114 5570 166
rect 7895 114 7947 166
rect 5326 104 5438 106
rect 5266 -10 5438 104
rect 5832 -2 6914 64
rect 5266 -108 5370 -10
rect 4918 -484 4994 -408
rect 5094 -722 5146 -670
rect 4746 -1300 4822 -1054
rect 4950 -1359 5027 -1282
rect 4732 -1602 4809 -1525
rect 4950 -1602 5027 -1525
rect 3026 -2232 3080 -2178
rect 948 -3290 1042 -3204
rect 1398 -3288 1492 -3202
rect 1856 -3290 1950 -3204
rect 2314 -3288 2408 -3202
rect 3942 -2244 4022 -2164
rect 4688 -2690 4798 -2614
rect 5094 -2678 5146 -2626
rect 5920 -1120 6052 -1068
rect 6178 -1120 6310 -1068
rect 6436 -1122 6568 -1070
rect 6694 -1130 6826 -1074
rect 7468 -1120 7600 -1064
rect 7726 -1120 7858 -1064
rect 7984 -1120 8116 -1064
rect 8242 -1120 8374 -1064
rect 9016 -1120 9148 -1064
rect 9274 -1120 9406 -1064
rect 9532 -1120 9664 -1064
rect 9790 -1120 9922 -1064
rect 10048 -1120 10180 -1064
rect 10965 1 11067 103
rect 10306 -1120 10438 -1064
rect 10564 -1120 10696 -1064
rect 10822 -1120 10954 -1064
rect 11080 -1120 11212 -1064
rect 11338 -1120 11470 -1064
rect 11596 -1120 11728 -1064
rect 11854 -1120 11986 -1064
rect 12112 -1120 12244 -1064
rect 12370 -1120 12502 -1064
rect 12628 -1120 12760 -1064
rect 13526 -830 13598 -758
rect 12886 -1120 13018 -1064
rect 6208 -1674 6260 -1622
rect 5290 -3146 5482 -3040
rect 2770 -3290 2864 -3204
rect -4132 -3510 -4080 -3458
rect 5320 -3510 5372 -3458
rect -4267 -3597 -4213 -3543
rect 6824 -1686 6890 -1614
rect 7340 -1686 7406 -1614
rect 7856 -1686 7922 -1614
rect 8888 -1686 8954 -1614
rect 9920 -1686 9986 -1614
rect 10952 -1686 11018 -1614
rect 13527 -1357 13598 -1286
rect 13788 2631 13843 2686
rect 15618 3332 15670 3384
rect 13920 2416 13972 2468
rect 14700 2416 14752 2468
rect 16576 2372 16628 2424
rect 18106 4520 18186 4600
rect 18760 4522 18884 4574
rect 19018 4522 19142 4574
rect 19276 4522 19400 4574
rect 19534 4522 19658 4574
rect 20308 3600 20432 3652
rect 20566 3600 20690 3652
rect 20824 3600 20948 3652
rect 21082 3600 21206 3652
rect 21853 3478 21932 3557
rect 18106 3034 18186 3114
rect 18923 3219 18981 3277
rect 17690 2372 17742 2424
rect 14524 2090 14652 2142
rect 14782 2090 14910 2142
rect 15040 2090 15168 2142
rect 15298 2090 15426 2142
rect 15556 2090 15684 2142
rect 15814 2090 15942 2142
rect 16588 2090 16718 2142
rect 16846 2090 16976 2142
rect 17102 2090 17232 2142
rect 16728 961 16802 1035
rect 17911 2355 17977 2421
rect 21702 3272 21774 3344
rect 17911 2081 17977 2147
rect 18624 2090 18748 2144
rect 17690 960 17742 1012
rect 19581 961 19655 1035
rect 15920 806 15992 878
rect 21580 806 21652 878
rect 13920 638 13972 690
rect 14524 -820 14648 -768
rect 15166 638 15218 690
rect 14782 -820 14906 -768
rect 15040 -820 15164 -768
rect 15298 -820 15422 -768
rect 15556 -820 15680 -768
rect 15814 -820 15938 -768
rect 16072 -820 16196 -768
rect 16330 -820 16454 -768
rect 16588 -820 16712 -768
rect 16846 -820 16970 -768
rect 17104 -820 17228 -768
rect 17362 -820 17486 -768
rect 18136 -820 18260 -768
rect 18394 -820 18518 -768
rect 18652 -820 18776 -768
rect 18910 -820 19034 -768
rect 19168 -820 19292 -768
rect 19426 -820 19550 -768
rect 19684 -820 19808 -768
rect 19942 -820 20066 -768
rect 20200 -820 20324 -768
rect 20458 -820 20582 -768
rect 20716 -820 20840 -768
rect 20974 -820 21098 -768
rect 13788 -1279 13843 -1224
rect 13982 -1270 14034 -1218
rect 14688 -1270 14742 -1218
rect 13660 -1438 13712 -1386
rect 11680 -1686 11882 -1618
rect 11984 -1686 12050 -1614
rect 12500 -1686 12566 -1614
rect 13016 -1686 13082 -1614
rect 8148 -1738 8406 -1734
rect 8148 -1790 8432 -1738
rect 8148 -1800 8406 -1790
rect 6920 -3124 9364 -3064
rect 9510 -3124 10396 -3064
rect 11474 -1786 11528 -1734
rect 10546 -3124 12986 -3064
rect 6326 -3250 6388 -3188
rect 9410 -3240 9464 -3188
rect 10442 -3240 10496 -3188
rect 13662 -3762 13714 -3710
rect 16236 -1270 16290 -1218
rect 16752 -1270 16806 -1218
rect 18300 -1270 18354 -1218
rect 18816 -1270 18870 -1218
rect 15204 -1436 15258 -1384
rect 15720 -1436 15774 -1384
rect 15924 -1450 16076 -1378
rect 17268 -1436 17322 -1384
rect 17784 -1436 17838 -1384
rect 19518 -1280 19698 -1208
rect 20364 -1270 20418 -1218
rect 19332 -1436 19386 -1384
rect 19846 -1436 19900 -1384
rect 22720 12146 22799 12225
rect 22584 11792 22656 11864
rect 22708 11304 22771 11367
rect 22402 9496 22454 9548
rect 22562 9376 22614 9428
rect 22402 8222 22454 8274
rect 22200 3478 22279 3557
rect 22030 3272 22102 3344
rect 22028 3034 22108 3114
rect 23339 11072 23400 11133
rect 23461 13841 23519 13899
rect 23589 13689 23655 13755
rect 23589 11683 23655 11749
rect 24136 11696 24260 11748
rect 24394 11696 24518 11748
rect 24652 11696 24776 11748
rect 25426 11696 25550 11748
rect 25684 11696 25808 11748
rect 25942 11696 26066 11748
rect 26200 11696 26324 11748
rect 26458 11696 26582 11748
rect 26716 11696 26840 11748
rect 26974 11696 27098 11748
rect 27232 11696 27356 11748
rect 26364 11514 26416 11566
rect 27490 11696 27614 11748
rect 27748 11696 28130 11748
rect 28264 11696 28646 11748
rect 28780 11696 29162 11748
rect 29296 11696 29420 11748
rect 29554 11696 29678 11748
rect 29812 11696 29936 11748
rect 26882 11514 26934 11566
rect 27397 11514 27449 11566
rect 27650 11516 27702 11568
rect 25332 11398 25384 11450
rect 25849 11398 25901 11450
rect 24302 11264 24354 11316
rect 24451 11264 24503 11316
rect 24817 11264 24869 11316
rect 23438 10924 23542 11004
rect 29464 11512 29516 11566
rect 30070 11696 30194 11748
rect 30328 11696 30452 11748
rect 30586 11696 30710 11748
rect 30844 11696 30968 11748
rect 29978 11512 30030 11564
rect 31102 11696 31226 11748
rect 31360 11696 31484 11748
rect 32134 11696 32258 11748
rect 32392 11696 32516 11748
rect 32650 11696 32774 11748
rect 30494 11512 30546 11564
rect 29611 11398 29663 11450
rect 31008 11396 31060 11450
rect 28428 11158 28480 11210
rect 31524 11396 31576 11448
rect 32042 11264 32094 11316
rect 32556 11264 32608 11316
rect 31676 11158 31728 11210
rect 29605 11006 29666 11067
rect 23254 9776 23378 9828
rect 23512 9776 23636 9828
rect 23770 9776 23894 9828
rect 24028 9776 24152 9828
rect 24286 9776 24410 9828
rect 24544 9776 24668 9828
rect 25318 9776 25442 9828
rect 25576 9776 25700 9828
rect 25834 9776 25958 9828
rect 26092 9776 26216 9828
rect 26350 9776 26474 9828
rect 26608 9776 26732 9828
rect 26866 9776 26990 9828
rect 27124 9776 27248 9828
rect 27382 9776 27506 9828
rect 27640 9776 27764 9828
rect 27898 9776 28022 9828
rect 28156 9776 28280 9828
rect 28930 9776 29054 9828
rect 29188 9776 29312 9828
rect 29446 9776 29570 9828
rect 29704 9776 29828 9828
rect 29962 9776 30086 9828
rect 30220 9776 30344 9828
rect 30994 9776 32410 9828
rect 26480 9496 26532 9548
rect 31920 9514 31996 9590
rect 33326 9514 33402 9590
rect 29624 9376 29676 9428
rect 23642 8712 23714 8784
rect 24252 8722 24376 8774
rect 24510 8722 24634 8774
rect 24768 8722 24892 8774
rect 25026 8722 25150 8774
rect 25284 8722 25408 8774
rect 25542 8722 25666 8774
rect 25800 8722 25924 8774
rect 26058 8722 26182 8774
rect 26316 8722 26440 8774
rect 26574 8722 26698 8774
rect 26832 8722 26956 8774
rect 27090 8722 27214 8774
rect 27348 8722 27472 8774
rect 27606 8722 27730 8774
rect 27864 8722 27988 8774
rect 28122 8722 28246 8774
rect 28380 8722 28504 8774
rect 28638 8722 28762 8774
rect 28896 8722 29020 8774
rect 29154 8722 29278 8774
rect 29412 8722 29536 8774
rect 29670 8722 29794 8774
rect 29928 8722 30052 8774
rect 30186 8722 30310 8774
rect 30444 8722 30568 8774
rect 30702 8722 30826 8774
rect 30960 8722 31084 8774
rect 31218 8722 31342 8774
rect 31476 8722 31600 8774
rect 31734 8722 31858 8774
rect 31992 8722 32116 8774
rect 32250 8722 32374 8774
rect 23376 8364 23428 8416
rect 22708 8097 22771 8160
rect 22707 4921 22777 4991
rect 23642 4752 23714 4824
rect 22555 2355 22621 2421
rect 28326 2666 28650 2948
rect 30842 2032 30902 2092
rect 22419 951 22505 1037
rect 22419 -426 22505 -340
rect 32006 2032 32066 2092
rect 32714 1910 32810 2006
rect 32854 1654 32950 1750
rect 22996 -416 31120 -350
rect 22028 -608 22108 -528
rect 21853 -756 21932 -677
rect 21702 -896 21774 -824
rect 14524 -2972 20582 -2920
rect 21580 -2982 21652 -2910
rect 14682 -3597 14737 -3542
rect 13982 -3876 14034 -3824
rect 6208 -3972 6260 -3920
rect 23822 -966 25936 -910
rect 26918 -966 29032 -910
rect 30014 -966 32128 -910
rect 22624 -1110 22748 -1058
rect 22882 -1110 23006 -1058
rect 22534 -1868 22600 -1796
rect 21871 -1946 21923 -1894
rect 21705 -4102 21778 -4029
rect 23656 -1110 23780 -1058
rect 23914 -1110 24038 -1058
rect 24172 -1110 24296 -1058
rect 24430 -1110 24554 -1058
rect 24688 -1110 24812 -1058
rect 24946 -1110 25070 -1058
rect 25204 -1110 25328 -1058
rect 25462 -1110 25586 -1058
rect 25718 -1110 25842 -1058
rect 25978 -1110 26102 -1058
rect 26752 -1110 26876 -1058
rect 27008 -1110 27132 -1058
rect 27268 -1110 27392 -1058
rect 27526 -1110 27650 -1058
rect 27784 -1110 27908 -1058
rect 28042 -1110 28166 -1058
rect 28300 -1110 28424 -1058
rect 28558 -1110 28682 -1058
rect 28816 -1110 28940 -1058
rect 29074 -1110 29198 -1058
rect 29848 -1110 29972 -1058
rect 23050 -1868 23116 -1796
rect 24598 -1950 24664 -1878
rect 23566 -2064 23632 -1992
rect 24082 -2064 24148 -1992
rect 30106 -1110 30230 -1058
rect 30364 -1110 30488 -1058
rect 30622 -1110 30746 -1058
rect 30880 -1110 31004 -1058
rect 31138 -1110 31262 -1058
rect 31396 -1110 31520 -1058
rect 31654 -1110 31778 -1058
rect 31912 -1110 32036 -1058
rect 33326 -976 33402 -900
rect 32170 -1110 32294 -1058
rect 25630 -1864 25696 -1792
rect 25114 -1950 25180 -1878
rect 24850 -2052 24908 -2000
rect 26146 -1950 26212 -1878
rect 28728 -1858 28792 -1796
rect 31040 -1848 31104 -1786
rect 31308 -1854 31368 -1792
rect 31824 -1854 31884 -1792
rect 27942 -1954 28010 -1898
rect 28210 -1964 28274 -1902
rect 26662 -2064 26728 -1992
rect 22634 -3006 22758 -2952
rect 22817 -3011 22875 -2953
rect 22892 -3006 23016 -2952
rect 23150 -3006 23274 -2952
rect 23408 -3006 23532 -2952
rect 23666 -3006 23790 -2952
rect 23924 -3006 24048 -2952
rect 24696 -3006 24820 -2952
rect 24956 -3006 25080 -2952
rect 25216 -3006 25340 -2952
rect 25474 -3006 25598 -2952
rect 25730 -3006 25854 -2952
rect 25988 -3006 26112 -2952
rect 27696 -2082 27760 -2020
rect 27174 -2164 27250 -2094
rect 26244 -3008 26368 -2954
rect 26506 -3008 26630 -2954
rect 26762 -3008 26886 -2954
rect 27022 -3008 27404 -2954
rect 27538 -3008 27662 -2954
rect 27794 -3008 27918 -2954
rect 29244 -1962 29304 -1900
rect 29760 -1960 29820 -1898
rect 30274 -2080 30338 -2018
rect 30792 -2080 30856 -2018
rect 28054 -3010 28178 -2956
rect 28310 -3008 28434 -2954
rect 28568 -3008 28692 -2954
rect 28826 -3008 28950 -2954
rect 29084 -3008 29208 -2954
rect 29342 -3008 29466 -2954
rect 29600 -3008 29724 -2954
rect 30374 -3006 30498 -2952
rect 30632 -3006 30756 -2952
rect 30890 -3006 31014 -2952
rect 31148 -3006 31272 -2952
rect 31406 -3006 31530 -2952
rect 31664 -3006 31788 -2952
rect 21870 -4267 21922 -4215
rect -5137 -4399 -5079 -4341
rect 22817 -4399 22875 -4341
<< metal2 >>
rect -4188 14039 -4182 14100
rect -4121 14039 23339 14100
rect 23400 14039 23406 14100
rect -3953 13841 -3947 13899
rect -3889 13841 23461 13899
rect 23519 13841 23525 13899
rect -5332 13786 -5248 13792
rect -5248 13702 -5190 13786
rect -5106 13702 -5097 13786
rect -5332 13696 -5248 13702
rect -3777 13689 -3771 13755
rect -3705 13689 23589 13755
rect 23655 13689 23661 13755
rect -3567 13473 -3561 13535
rect -3499 13473 17467 13535
rect 17529 13473 17535 13535
rect -3451 13341 -3445 13399
rect -3387 13341 17191 13399
rect 17249 13341 17255 13399
rect -3340 13198 -3334 13266
rect -3266 13265 -2772 13266
rect -3266 13199 16971 13265
rect 17037 13199 17043 13265
rect -3266 13198 -2772 13199
rect -3214 13074 -3208 13134
rect -3148 13074 12756 13134
rect 12696 13018 12756 13074
rect 2776 12928 2782 12980
rect 2834 12979 2840 12980
rect 11548 12979 11554 12980
rect 2834 12929 11554 12979
rect 2834 12928 2840 12929
rect 11548 12928 11554 12929
rect 11606 12928 11612 12980
rect 11802 12942 11808 13014
rect 11880 12942 12478 13014
rect 12550 12942 12559 13014
rect 12688 12946 12694 13018
rect 12766 13013 13418 13018
rect 12766 12951 13351 13013
rect 13413 12951 13422 13013
rect 12766 12946 13418 12951
rect 12696 12936 12756 12946
rect 14159 12943 14211 12945
rect 14675 12943 14727 12944
rect 14158 12935 20151 12943
rect 14158 12883 14159 12935
rect 14211 12934 20151 12935
rect 14211 12883 14675 12934
rect 14158 12882 14675 12883
rect 14727 12933 20151 12934
rect 14727 12882 15707 12933
rect 14158 12881 15707 12882
rect 15759 12881 16223 12933
rect 16275 12929 20151 12933
rect 16275 12881 17191 12929
rect 14158 12873 17191 12881
rect 14675 12872 14727 12873
rect 15707 12871 15759 12873
rect 16223 12871 16275 12873
rect 17185 12871 17191 12873
rect 17249 12873 20151 12929
rect 20221 12873 20227 12943
rect 17249 12871 17255 12873
rect -2922 12772 -2916 12832
rect -2856 12772 2186 12832
rect 2246 12772 2252 12832
rect 13337 12729 13346 12801
rect 13418 12791 18348 12801
rect 13418 12739 15191 12791
rect 15243 12739 18348 12791
rect 13418 12729 18348 12739
rect 18420 12729 18426 12801
rect 9516 12642 9576 12648
rect -3086 12560 -3080 12632
rect -3008 12622 1670 12632
rect -3008 12570 -2324 12622
rect -2200 12570 -2066 12622
rect -1942 12570 -1808 12622
rect -1684 12570 -1550 12622
rect -1426 12570 -1292 12622
rect -1168 12570 -1034 12622
rect -910 12570 -776 12622
rect -652 12570 -518 12622
rect -394 12570 -260 12622
rect -136 12570 -2 12622
rect 122 12570 256 12622
rect 380 12570 514 12622
rect 638 12570 772 12622
rect 896 12570 1030 12622
rect 1154 12570 1288 12622
rect 1412 12570 1546 12622
rect 2180 12582 2186 12642
rect 2246 12582 9516 12642
rect 9516 12576 9576 12582
rect -3008 12560 1670 12570
rect 2590 12436 2596 12516
rect 2676 12498 8422 12516
rect 2676 12446 3396 12498
rect 3520 12446 3654 12498
rect 3778 12446 3912 12498
rect 4036 12446 4170 12498
rect 4294 12446 4428 12498
rect 4552 12446 4686 12498
rect 4810 12446 4944 12498
rect 5068 12446 5202 12498
rect 5326 12446 5460 12498
rect 5584 12446 5718 12498
rect 5842 12446 5976 12498
rect 6100 12446 6234 12498
rect 6358 12446 6492 12498
rect 6616 12446 6750 12498
rect 6874 12446 7008 12498
rect 7132 12446 7266 12498
rect 7390 12446 7524 12498
rect 7648 12446 7782 12498
rect 7906 12446 8040 12498
rect 8164 12446 8298 12498
rect 2676 12436 8422 12446
rect 9748 12500 11808 12510
rect 9800 12448 9914 12500
rect 10112 12448 10230 12500
rect 10428 12448 10546 12500
rect 10744 12448 10862 12500
rect 10914 12448 11808 12500
rect 9748 12438 11808 12448
rect 11880 12438 11886 12510
rect 22376 12225 22385 12235
rect 12308 12156 12398 12166
rect 22194 12146 22200 12225
rect 22279 12153 22385 12225
rect 22467 12225 22476 12235
rect 22467 12153 22720 12225
rect 22279 12146 22720 12153
rect 22799 12146 22805 12225
rect 12412 12115 21152 12118
rect 12412 12049 16971 12115
rect 17037 12108 21152 12115
rect 17037 12056 18190 12108
rect 18314 12056 18448 12108
rect 18572 12056 19222 12108
rect 19346 12056 19480 12108
rect 19604 12056 19738 12108
rect 19862 12056 19996 12108
rect 20120 12056 20254 12108
rect 20378 12056 20512 12108
rect 20636 12056 20770 12108
rect 20894 12056 21028 12108
rect 17037 12049 21152 12056
rect 12412 12046 21152 12049
rect 12308 12000 12398 12010
rect 12152 11850 12260 11860
rect 13380 11859 22584 11864
rect 12976 11850 13084 11858
rect 11321 11762 11330 11850
rect 11418 11768 12152 11850
rect 12260 11848 13084 11850
rect 12260 11768 12976 11848
rect 11418 11766 12976 11768
rect 13376 11797 13385 11859
rect 13447 11797 22584 11859
rect 13380 11792 22584 11797
rect 22656 11792 22662 11864
rect 11418 11762 13084 11766
rect 12152 11758 12260 11762
rect 12976 11756 13084 11762
rect 24136 11749 32774 11758
rect 23583 11683 23589 11749
rect 23655 11748 32774 11749
rect 23655 11696 24136 11748
rect 24260 11696 24394 11748
rect 24518 11696 24652 11748
rect 24776 11696 25426 11748
rect 25550 11696 25684 11748
rect 25808 11696 25942 11748
rect 26066 11696 26200 11748
rect 26324 11696 26458 11748
rect 26582 11696 26716 11748
rect 26840 11696 26974 11748
rect 27098 11696 27232 11748
rect 27356 11696 27490 11748
rect 27614 11696 27748 11748
rect 28130 11696 28264 11748
rect 28646 11696 28780 11748
rect 29162 11696 29296 11748
rect 29420 11696 29554 11748
rect 29678 11696 29812 11748
rect 29936 11696 30070 11748
rect 30194 11696 30328 11748
rect 30452 11696 30586 11748
rect 30710 11696 30844 11748
rect 30968 11696 31102 11748
rect 31226 11696 31360 11748
rect 31484 11696 32134 11748
rect 32258 11696 32392 11748
rect 32516 11696 32650 11748
rect 23655 11686 32774 11696
rect 23655 11683 24311 11686
rect 27397 11566 27449 11572
rect 11810 11556 11926 11566
rect 11554 11546 11606 11552
rect 11606 11495 11810 11545
rect 11554 11488 11606 11494
rect 18346 11545 18352 11546
rect 11926 11539 18352 11545
rect 11926 11495 17467 11539
rect 11810 11476 11926 11486
rect 17461 11477 17467 11495
rect 17529 11495 18352 11539
rect 17529 11477 17535 11495
rect 18346 11494 18352 11495
rect 18404 11494 18410 11546
rect 26358 11514 26364 11566
rect 26416 11563 26422 11566
rect 26876 11563 26882 11566
rect 26416 11517 26882 11563
rect 26416 11514 26422 11517
rect 26876 11514 26882 11517
rect 26934 11563 26940 11566
rect 26934 11517 27397 11563
rect 26934 11514 26940 11517
rect 27644 11563 27650 11568
rect 27449 11517 27650 11563
rect 27644 11516 27650 11517
rect 27702 11563 27708 11568
rect 29458 11563 29464 11566
rect 27702 11517 29464 11563
rect 27702 11516 27708 11517
rect 27397 11508 27449 11514
rect 29458 11512 29464 11517
rect 29516 11561 29522 11566
rect 29972 11561 29978 11564
rect 29516 11515 29978 11561
rect 29516 11512 29522 11515
rect 29972 11512 29978 11515
rect 30030 11561 30036 11564
rect 30488 11561 30494 11564
rect 30030 11515 30494 11561
rect 30030 11512 30036 11515
rect 30488 11512 30494 11515
rect 30546 11512 30552 11564
rect 11678 11328 11684 11400
rect 11756 11393 13380 11400
rect 11756 11331 12483 11393
rect 12545 11331 13380 11393
rect 11756 11328 13380 11331
rect 13452 11328 13461 11400
rect 25326 11398 25332 11450
rect 25384 11447 25390 11450
rect 25843 11447 25849 11450
rect 25384 11401 25849 11447
rect 25384 11398 25390 11401
rect 25843 11398 25849 11401
rect 25901 11447 25907 11450
rect 29605 11447 29611 11450
rect 25901 11401 29611 11447
rect 25901 11398 25907 11401
rect 29605 11398 29611 11401
rect 29663 11447 29669 11450
rect 31002 11447 31008 11450
rect 29663 11401 31008 11447
rect 29663 11398 29669 11401
rect 31002 11396 31008 11401
rect 31060 11445 31066 11450
rect 31518 11445 31524 11448
rect 31060 11399 31524 11445
rect 31060 11396 31066 11399
rect 31518 11396 31524 11399
rect 31576 11396 31582 11448
rect 19947 11304 19953 11367
rect 20016 11304 22708 11367
rect 22771 11304 22777 11367
rect 24296 11264 24302 11316
rect 24354 11313 24360 11316
rect 24445 11313 24451 11316
rect 24354 11267 24451 11313
rect 24354 11264 24360 11267
rect 24445 11264 24451 11267
rect 24503 11313 24509 11316
rect 24811 11313 24817 11316
rect 24503 11267 24817 11313
rect 24503 11264 24509 11267
rect 24811 11264 24817 11267
rect 24869 11313 24875 11316
rect 32036 11313 32042 11316
rect 24869 11267 32042 11313
rect 24869 11264 24875 11267
rect 32036 11264 32042 11267
rect 32094 11313 32100 11316
rect 32550 11313 32556 11316
rect 32094 11267 32556 11313
rect 32094 11264 32100 11267
rect 32550 11264 32556 11267
rect 32608 11264 32614 11316
rect 11544 11158 11550 11230
rect 11622 11220 21468 11230
rect 11622 11168 12314 11220
rect 12438 11168 12572 11220
rect 12696 11168 12830 11220
rect 12954 11168 13088 11220
rect 13212 11168 13346 11220
rect 13470 11168 13604 11220
rect 13728 11168 13862 11220
rect 13986 11168 14120 11220
rect 14244 11168 14378 11220
rect 14502 11168 14636 11220
rect 14760 11168 14894 11220
rect 15018 11168 15152 11220
rect 15276 11168 15410 11220
rect 15534 11168 15668 11220
rect 15792 11168 15926 11220
rect 16050 11168 16184 11220
rect 16308 11168 16442 11220
rect 16566 11168 16700 11220
rect 16824 11168 16958 11220
rect 17082 11168 17216 11220
rect 17340 11168 17474 11220
rect 17598 11168 17732 11220
rect 17856 11168 17990 11220
rect 18114 11168 18248 11220
rect 18372 11168 18506 11220
rect 18630 11168 18764 11220
rect 18888 11168 19022 11220
rect 19146 11168 19280 11220
rect 19404 11168 19538 11220
rect 19662 11168 19796 11220
rect 19920 11168 20054 11220
rect 20178 11168 20312 11220
rect 20436 11168 20570 11220
rect 20694 11168 20828 11220
rect 20952 11168 21086 11220
rect 21210 11168 21344 11220
rect 11622 11158 21468 11168
rect 28422 11158 28428 11210
rect 28480 11208 28486 11210
rect 31670 11208 31676 11210
rect 28480 11160 31676 11208
rect 28480 11158 28486 11160
rect 31670 11158 31676 11160
rect 31728 11158 31734 11210
rect 23333 11072 23339 11133
rect 23400 11072 28328 11133
rect 28267 11067 28328 11072
rect 29588 11067 29686 11080
rect 23438 11004 23542 11014
rect 28267 11006 29605 11067
rect 29666 11006 29686 11067
rect 29588 10990 29686 11006
rect 23438 10914 23542 10924
rect 2699 10309 3777 10311
rect 6882 10309 6888 10310
rect 2699 10308 3560 10309
rect 2693 10252 2702 10308
rect 2758 10255 3560 10308
rect 3614 10307 4592 10309
rect 3614 10255 4076 10307
rect 2758 10252 3777 10255
rect 4070 10253 4076 10255
rect 4130 10255 4592 10307
rect 4646 10255 5108 10309
rect 5162 10307 6888 10309
rect 5162 10255 6656 10307
rect 4130 10253 4136 10255
rect 6650 10253 6656 10255
rect 6710 10258 6888 10307
rect 6940 10309 6946 10310
rect 6940 10258 7172 10309
rect 6710 10255 7172 10258
rect 7226 10255 7688 10309
rect 7742 10255 8203 10309
rect 8257 10255 8263 10309
rect 6710 10253 6716 10255
rect 2699 10249 3777 10252
rect 3793 10147 3799 10201
rect 3853 10147 5883 10201
rect 5937 10147 5943 10201
rect 2412 9880 2418 9932
rect 2470 9931 2476 9932
rect 9764 9931 9770 9932
rect 2470 9881 9770 9931
rect 2470 9880 2476 9881
rect 9764 9880 9770 9881
rect 9822 9880 9828 9932
rect 23461 9838 23519 10914
rect 23254 9828 32410 9838
rect 2250 9750 2256 9802
rect 2308 9801 2314 9802
rect 9548 9801 9554 9802
rect 2308 9751 9554 9801
rect 2308 9750 2314 9751
rect 9548 9750 9554 9751
rect 9606 9750 9612 9802
rect 23378 9776 23512 9828
rect 23636 9776 23770 9828
rect 23894 9776 24028 9828
rect 24152 9776 24286 9828
rect 24410 9776 24544 9828
rect 24668 9776 25318 9828
rect 25442 9776 25576 9828
rect 25700 9776 25834 9828
rect 25958 9776 26092 9828
rect 26216 9776 26350 9828
rect 26474 9776 26608 9828
rect 26732 9776 26866 9828
rect 26990 9776 27124 9828
rect 27248 9776 27382 9828
rect 27506 9776 27640 9828
rect 27764 9776 27898 9828
rect 28022 9776 28156 9828
rect 28280 9776 28930 9828
rect 29054 9776 29188 9828
rect 29312 9776 29446 9828
rect 29570 9776 29704 9828
rect 29828 9776 29962 9828
rect 30086 9776 30220 9828
rect 30344 9776 30994 9828
rect 23254 9766 32410 9776
rect 23461 9757 23519 9766
rect 3384 9541 11684 9548
rect 2508 9538 11684 9541
rect 2502 9482 2511 9538
rect 2567 9486 3384 9538
rect 3508 9486 3642 9538
rect 3766 9486 3900 9538
rect 4024 9486 4158 9538
rect 4282 9486 4932 9538
rect 5056 9486 5190 9538
rect 5314 9486 5448 9538
rect 5572 9486 5706 9538
rect 5830 9486 5964 9538
rect 6088 9486 6222 9538
rect 6346 9486 6480 9538
rect 6604 9486 6738 9538
rect 6862 9486 6996 9538
rect 7120 9486 7254 9538
rect 7378 9486 7512 9538
rect 7636 9486 7770 9538
rect 7894 9486 8028 9538
rect 8152 9486 8286 9538
rect 8410 9486 8544 9538
rect 8668 9486 8802 9538
rect 8926 9486 11684 9538
rect 2567 9482 11684 9486
rect 2508 9479 11684 9482
rect 3384 9476 11684 9479
rect 11756 9476 11762 9548
rect 22396 9496 22402 9548
rect 22454 9547 22460 9548
rect 26474 9547 26480 9548
rect 22454 9497 26480 9547
rect 22454 9496 22460 9497
rect 26474 9496 26480 9497
rect 26532 9496 26538 9548
rect 31914 9514 31920 9590
rect 31996 9514 33326 9590
rect 33402 9514 33408 9590
rect 22556 9376 22562 9428
rect 22614 9427 22620 9428
rect 29618 9427 29624 9428
rect 22614 9377 29624 9427
rect 22614 9376 22620 9377
rect 29618 9376 29624 9377
rect 29676 9376 29682 9428
rect -992 8974 -986 8976
rect -3086 8902 -3080 8974
rect -3008 8920 -986 8974
rect -930 8974 -924 8976
rect -930 8920 1894 8974
rect -3008 8902 1894 8920
rect 1966 8902 1972 8974
rect 30573 8874 30582 8970
rect 30678 8965 33522 8970
rect 30678 8879 33431 8965
rect 33517 8879 33526 8965
rect 30678 8874 33522 8879
rect -2919 8755 -2913 8809
rect -2859 8755 1689 8809
rect 1743 8755 1749 8809
rect 23642 8784 23714 8790
rect 30578 8784 30587 8793
rect 23714 8774 30587 8784
rect 23714 8722 24252 8774
rect 24376 8722 24510 8774
rect 24634 8722 24768 8774
rect 24892 8722 25026 8774
rect 25150 8722 25284 8774
rect 25408 8722 25542 8774
rect 25666 8722 25800 8774
rect 25924 8722 26058 8774
rect 26182 8722 26316 8774
rect 26440 8722 26574 8774
rect 26698 8722 26832 8774
rect 26956 8722 27090 8774
rect 27214 8722 27348 8774
rect 27472 8722 27606 8774
rect 27730 8722 27864 8774
rect 27988 8722 28122 8774
rect 28246 8722 28380 8774
rect 28504 8722 28638 8774
rect 28762 8722 28896 8774
rect 29020 8722 29154 8774
rect 29278 8722 29412 8774
rect 29536 8722 29670 8774
rect 29794 8722 29928 8774
rect 30052 8722 30186 8774
rect 30310 8722 30444 8774
rect 30568 8722 30587 8774
rect 23714 8712 30587 8722
rect 23642 8706 23714 8712
rect 30578 8707 30587 8712
rect 30673 8784 30682 8793
rect 30673 8774 32374 8784
rect 30673 8722 30702 8774
rect 30826 8722 30960 8774
rect 31084 8722 31218 8774
rect 31342 8722 31476 8774
rect 31600 8722 31734 8774
rect 31858 8722 31992 8774
rect 32116 8722 32250 8774
rect 30673 8712 32374 8722
rect 30673 8707 30682 8712
rect -3214 8646 -3208 8706
rect -3148 8646 322 8706
rect 382 8646 388 8706
rect 427 8606 433 8607
rect -3340 8538 -3334 8606
rect -3266 8538 433 8606
rect 427 8537 433 8538
rect 503 8537 509 8607
rect -3451 8435 -3445 8493
rect -3387 8435 -533 8493
rect -475 8435 -469 8493
rect 785 8479 791 8541
rect 853 8479 2699 8541
rect 2761 8479 2770 8541
rect 10892 8512 10898 8591
rect 10977 8512 13666 8591
rect 13745 8512 13751 8591
rect -3567 8317 -3561 8379
rect -3499 8317 -653 8379
rect -591 8317 -585 8379
rect 2084 8356 2090 8432
rect 2166 8356 2780 8432
rect 2856 8356 2862 8432
rect 9548 8364 9554 8416
rect 9606 8415 9612 8416
rect 23370 8415 23376 8416
rect 9606 8365 23376 8415
rect 9606 8364 9612 8365
rect 23370 8364 23376 8365
rect 23428 8364 23434 8416
rect 9764 8222 9770 8274
rect 9822 8273 9828 8274
rect 22396 8273 22402 8274
rect 9822 8223 22402 8273
rect 9822 8222 9828 8223
rect 22396 8222 22402 8223
rect 22454 8222 22460 8274
rect -3771 8131 -3705 8137
rect -3705 8065 -1607 8131
rect -1541 8065 -1535 8131
rect 18677 8097 18683 8160
rect 18746 8097 22708 8160
rect 22771 8097 22777 8160
rect -3771 8059 -3705 8065
rect 11178 8010 11184 8082
rect 11256 8010 11550 8082
rect 11622 8010 11628 8082
rect 11814 7938 22380 7960
rect -3953 7851 -3947 7909
rect -3889 7851 -1755 7909
rect -1697 7851 -1691 7909
rect 11938 7886 12072 7938
rect 12196 7886 12330 7938
rect 12454 7886 12588 7938
rect 12712 7886 12846 7938
rect 12970 7886 13104 7938
rect 13228 7886 13362 7938
rect 13486 7886 13620 7938
rect 13744 7886 13878 7938
rect 14002 7886 14136 7938
rect 14260 7886 14394 7938
rect 14518 7886 14652 7938
rect 14776 7886 14910 7938
rect 15034 7886 15168 7938
rect 15292 7886 15426 7938
rect 15550 7886 15684 7938
rect 15808 7886 15942 7938
rect 16066 7886 16200 7938
rect 16324 7886 16974 7938
rect 17098 7886 17232 7938
rect 17356 7886 17490 7938
rect 17614 7886 17748 7938
rect 17872 7886 18006 7938
rect 18130 7886 18264 7938
rect 18388 7886 18522 7938
rect 18646 7886 18780 7938
rect 18904 7886 19038 7938
rect 19162 7886 19296 7938
rect 19420 7886 19554 7938
rect 19678 7886 19812 7938
rect 19936 7886 20070 7938
rect 20194 7886 20328 7938
rect 20452 7886 20586 7938
rect 20710 7886 20844 7938
rect 20968 7886 21102 7938
rect 21226 7886 21360 7938
rect 21484 7886 22380 7938
rect 11814 7868 22380 7886
rect 22472 7868 22481 7960
rect -4188 7633 -4182 7694
rect -4121 7633 -1918 7694
rect -1857 7633 -1851 7694
rect 2630 7428 2636 7480
rect 2688 7479 2694 7480
rect 3806 7479 3812 7480
rect 2688 7429 3812 7479
rect 2688 7428 2694 7429
rect 3806 7428 3812 7429
rect 3864 7428 3870 7480
rect 6596 7457 6602 7504
rect 6559 7388 6602 7457
rect 6718 7499 10026 7504
rect 6718 7393 9915 7499
rect 10021 7463 10030 7499
rect 10021 7401 10213 7463
rect 10275 7401 10281 7463
rect 10021 7393 10030 7401
rect 6718 7388 10026 7393
rect 6559 7387 6985 7388
rect -4386 7174 -3900 7310
rect 1435 7293 1441 7387
rect 1535 7293 6985 7387
rect 2332 7206 10280 7210
rect -3775 7174 -3709 7178
rect -4386 7169 -3704 7174
rect -4386 7103 -3775 7169
rect -3709 7103 -3704 7169
rect 2327 7150 2336 7206
rect 2392 7150 10280 7206
rect 2332 7146 10280 7150
rect 10344 7146 10350 7210
rect -4386 7098 -3704 7103
rect -4386 6810 -3900 7098
rect -3775 7094 -3709 7098
rect -1613 7009 -1607 7075
rect -1541 7009 -913 7075
rect -847 7009 -841 7075
rect 790 7007 796 7068
rect 857 7007 2509 7068
rect 2570 7007 2579 7068
rect 2827 6996 2836 7052
rect 2892 7051 2901 7052
rect 2892 6997 10915 7051
rect 10969 6997 10975 7051
rect 2892 6996 2901 6997
rect 3338 6954 11034 6956
rect 3338 6904 10138 6954
rect -1761 6837 -1755 6895
rect -1697 6837 -1581 6895
rect -1523 6837 -1517 6895
rect 2524 6884 2834 6886
rect 2517 6828 2526 6884
rect 2582 6828 2834 6884
rect 2524 6826 2834 6828
rect 2894 6826 2903 6886
rect -4392 6294 -3906 6700
rect 3254 6616 3310 6626
rect -3818 6294 -3812 6308
rect -4392 6244 -3812 6294
rect -3748 6294 -3742 6308
rect -3328 6294 -3272 6301
rect -3748 6292 -3270 6294
rect -3748 6244 -3328 6292
rect -4392 6236 -3328 6244
rect -3272 6236 -3270 6292
rect -4392 6234 -3270 6236
rect -4392 6200 -3906 6234
rect -3328 6227 -3272 6234
rect -1918 6095 -1857 6101
rect -4392 5592 -3906 6092
rect -1922 6034 -1918 6095
rect -1857 6094 -1699 6095
rect -1857 6034 -1760 6094
rect -1700 6034 -1694 6094
rect -1918 6028 -1857 6034
rect -3162 5964 -3076 5974
rect -3162 5890 -3076 5900
rect -2198 5958 -2140 5968
rect -3154 5846 -3090 5890
rect -2198 5882 -2140 5892
rect -2196 5846 -2142 5882
rect 2618 5876 2698 5886
rect -595 5867 -537 5873
rect -3154 5836 -2142 5846
rect -3154 5778 -2922 5836
rect -2374 5778 -2142 5836
rect -1587 5809 -1581 5867
rect -1523 5809 -595 5867
rect 792 5865 2618 5866
rect -595 5803 -537 5809
rect 787 5807 793 5865
rect 851 5807 2618 5865
rect 792 5806 2618 5807
rect 2618 5782 2698 5792
rect -3154 5770 -2142 5778
rect -3154 5768 -3090 5770
rect -2922 5768 -2142 5770
rect -2196 5766 -2142 5768
rect -4116 5550 -4056 5592
rect -4123 5494 -4114 5550
rect -4058 5494 -4049 5550
rect -4116 5492 -4056 5494
rect 3254 5384 3310 5394
rect 3512 6616 3568 6904
rect 3512 5336 3568 5394
rect 3770 6616 3826 6626
rect 3770 5384 3826 5394
rect 4028 6616 4084 6674
rect 4028 5234 4084 5394
rect 4286 6616 4342 6626
rect 4286 5384 4342 5394
rect 4544 6616 4600 6674
rect 4544 5234 4600 5394
rect 4802 6616 4858 6626
rect 4802 5384 4858 5394
rect 5060 6616 5116 6904
rect 5060 5336 5116 5394
rect 5318 6616 5374 6626
rect 5318 5384 5374 5394
rect 5576 6616 5632 6904
rect 5576 5336 5632 5394
rect 5834 6616 5890 6626
rect 5834 5384 5890 5394
rect 6092 6616 6148 6674
rect 6092 5234 6148 5394
rect 6350 6616 6406 6626
rect 6350 5384 6406 5394
rect 6608 6616 6664 6674
rect 6608 5234 6664 5394
rect 6866 6616 6922 6626
rect 6866 5384 6922 5394
rect 7124 6616 7180 6904
rect 7124 5336 7180 5394
rect 7382 6616 7438 6626
rect 7382 5384 7438 5394
rect 7640 6616 7696 6904
rect 7640 5336 7696 5394
rect 7898 6616 7954 6626
rect 7898 5384 7954 5394
rect 8156 6616 8212 6674
rect 8156 5234 8212 5394
rect 8414 6616 8470 6626
rect 8414 5384 8470 5394
rect 8672 6616 8728 6674
rect 8672 5234 8728 5394
rect 8930 6616 8986 6626
rect 8930 5384 8986 5394
rect 9188 6616 9244 6904
rect 10132 6902 10138 6904
rect 10190 6904 11034 6954
rect 11086 6904 11092 6956
rect 10190 6902 10196 6904
rect 9188 5336 9244 5394
rect 9446 6616 9502 6626
rect 9446 5384 9502 5394
rect 2980 5176 10449 5234
rect 10507 5176 10513 5234
rect 11178 5216 11184 5288
rect 11256 5216 14288 5288
rect 14360 5216 14366 5288
rect -5620 5022 -5614 5086
rect -5550 5022 -3812 5086
rect -3748 5022 -3742 5086
rect 3254 5012 3310 5022
rect -986 4942 -926 4948
rect -2514 4914 -2464 4918
rect -2274 4914 -2042 4922
rect -3254 4912 -2042 4914
rect -3254 4904 -2274 4912
rect -3022 4846 -2274 4904
rect -3022 4838 -2042 4846
rect -3254 4836 -2042 4838
rect -3254 4828 -3022 4836
rect -2832 4738 -2782 4836
rect -2514 4738 -2464 4836
rect -2844 4728 -2768 4738
rect -4332 4651 -3780 4656
rect -4336 4585 -4327 4651
rect -4261 4585 -3780 4651
rect -4332 4580 -3780 4585
rect -3704 4580 -3695 4656
rect -2844 4654 -2768 4664
rect -2528 4728 -2452 4738
rect -2528 4654 -2452 4664
rect -986 4660 -926 4882
rect 2515 4668 2524 4670
rect -1766 4600 -1760 4660
rect -1700 4600 -926 4660
rect 800 4612 806 4668
rect 862 4612 2524 4668
rect 2515 4610 2524 4612
rect 2584 4610 2593 4670
rect -8186 4249 -8122 4255
rect -6598 4249 -4028 4252
rect -8122 4188 -4028 4249
rect -3964 4188 -3958 4252
rect -8122 4185 -6569 4188
rect -8186 4179 -8122 4185
rect 3254 3780 3310 3790
rect 3512 5012 3568 5176
rect 3512 3732 3568 3790
rect 3770 5012 3826 5022
rect 3770 3780 3826 3790
rect 4028 5012 4084 5070
rect 4028 3534 4084 3790
rect 4286 5012 4342 5022
rect 4286 3780 4342 3790
rect 4544 5012 4600 5070
rect 4544 3534 4600 3790
rect 4802 5012 4858 5022
rect 4802 3780 4858 3790
rect 5060 5012 5116 5176
rect 5060 3732 5116 3790
rect 5318 5012 5374 5022
rect 5318 3780 5374 3790
rect 5576 5012 5632 5176
rect 5576 3732 5632 3790
rect 5834 5012 5890 5022
rect 5834 3780 5890 3790
rect 6092 5012 6148 5070
rect 6092 3534 6148 3790
rect 6350 5012 6406 5022
rect 6350 3780 6406 3790
rect 6608 5012 6664 5070
rect 6608 3534 6664 3790
rect 6866 5012 6922 5022
rect 6866 3780 6922 3790
rect 7124 5012 7180 5176
rect 7124 3732 7180 3790
rect 7382 5012 7438 5022
rect 7382 3780 7438 3790
rect 7640 5012 7696 5176
rect 7640 3732 7696 3790
rect 7898 5012 7954 5022
rect 7898 3780 7954 3790
rect 8156 5012 8212 5070
rect 8156 3534 8212 3790
rect 8414 5012 8470 5022
rect 8414 3780 8470 3790
rect 8672 5012 8728 5070
rect 8672 3534 8728 3790
rect 8930 5012 8986 5022
rect 8930 3780 8986 3790
rect 9188 5012 9244 5176
rect 11033 5118 13144 5120
rect 11028 5066 11034 5118
rect 11086 5066 13144 5118
rect 11033 5065 13144 5066
rect 13199 5065 13205 5120
rect 9188 3732 9244 3790
rect 9446 5012 9502 5022
rect 10274 4982 10350 4988
rect 12753 4982 12759 4991
rect 10274 4918 10280 4982
rect 10344 4921 12759 4982
rect 12829 4921 22707 4991
rect 22777 4921 22783 4991
rect 10344 4918 12870 4921
rect 10274 4910 10350 4918
rect 12554 4764 12560 4816
rect 12612 4814 12618 4816
rect 16186 4814 16192 4824
rect 12612 4772 16192 4814
rect 16244 4823 16250 4824
rect 17264 4823 17270 4828
rect 16244 4776 17270 4823
rect 17322 4823 17328 4828
rect 19186 4823 19200 4824
rect 17322 4776 19200 4823
rect 16244 4773 19200 4776
rect 16244 4772 16432 4773
rect 12612 4766 16432 4772
rect 19186 4772 19200 4773
rect 19252 4772 23642 4824
rect 12612 4764 12618 4766
rect 19186 4752 23642 4772
rect 23714 4752 23720 4824
rect 18100 4588 18106 4600
rect 13972 4585 18106 4588
rect 12409 4519 12415 4585
rect 12481 4578 18106 4585
rect 12481 4526 13972 4578
rect 14096 4526 14230 4578
rect 14354 4526 14488 4578
rect 14612 4526 14746 4578
rect 14870 4526 15004 4578
rect 15128 4526 15262 4578
rect 15386 4526 16036 4578
rect 16160 4526 16294 4578
rect 16418 4526 16552 4578
rect 16676 4526 18106 4578
rect 12481 4520 18106 4526
rect 18186 4588 18192 4600
rect 18186 4584 18890 4588
rect 18186 4574 19658 4584
rect 18186 4522 18760 4574
rect 18884 4522 19018 4574
rect 19142 4522 19276 4574
rect 19400 4522 19534 4574
rect 18186 4520 19658 4522
rect 12481 4519 19658 4520
rect 13972 4516 19658 4519
rect 18758 4512 19658 4516
rect 9446 3780 9502 3790
rect 20308 3652 21206 3662
rect 20432 3600 20566 3652
rect 20690 3600 20824 3652
rect 20948 3600 21082 3652
rect 20308 3590 21206 3600
rect 10443 3534 10449 3535
rect 358 3458 364 3522
rect 428 3458 2332 3522
rect 2396 3458 2405 3522
rect 3346 3482 10138 3534
rect 10190 3482 10202 3534
rect 10430 3482 10449 3534
rect 10443 3477 10449 3482
rect 10507 3534 10513 3535
rect 10507 3482 12994 3534
rect 13046 3482 13052 3534
rect 10507 3477 10513 3482
rect 21847 3478 21853 3557
rect 21932 3478 22200 3557
rect 22279 3478 22285 3557
rect 6041 3425 6120 3431
rect -4464 3349 -4210 3354
rect -6598 3346 -4210 3349
rect -8909 3284 -8903 3346
rect -8841 3287 -4210 3346
rect -8841 3284 -6443 3287
rect -4464 3282 -4210 3287
rect -4138 3282 -4132 3354
rect 6120 3346 10898 3425
rect 10977 3346 10983 3425
rect 6041 3340 6120 3346
rect 13310 3332 13316 3384
rect 13368 3332 15618 3384
rect 15670 3332 15676 3384
rect -1636 3324 -1580 3330
rect -1580 3268 -1234 3324
rect -1178 3268 -334 3324
rect -278 3268 94 3324
rect 150 3268 1056 3324
rect 1112 3268 1118 3324
rect -1636 3262 -1580 3268
rect 1519 3219 1525 3277
rect 1583 3219 18923 3277
rect 18981 3219 18987 3277
rect 21696 3272 21702 3344
rect 21774 3272 22030 3344
rect 22102 3272 22108 3344
rect -598 3110 -592 3162
rect -540 3160 -534 3162
rect 12554 3160 12560 3162
rect -540 3112 12560 3160
rect -540 3110 -534 3112
rect 12554 3110 12560 3112
rect 12612 3110 12618 3162
rect -4568 2996 -4562 3068
rect -4490 3060 -4010 3068
rect -4490 3000 -4116 3060
rect -4056 3054 -4010 3060
rect 4690 3058 13722 3060
rect 2828 3054 2834 3056
rect -4056 3006 2834 3054
rect -4056 3000 -4010 3006
rect 2828 3004 2834 3006
rect 2886 3054 2892 3056
rect 4690 3054 13664 3058
rect 2886 3006 13664 3054
rect 2886 3004 2892 3006
rect 4690 3002 13664 3006
rect 13720 3002 13729 3058
rect 18100 3034 18106 3114
rect 18186 3034 22028 3114
rect 22108 3034 22114 3114
rect 4690 3000 13722 3002
rect -4490 2996 -4010 3000
rect -1698 2964 -1644 2968
rect -3722 2962 -1631 2964
rect -3729 2906 -3720 2962
rect -3664 2958 -1631 2962
rect -3664 2906 -1698 2958
rect -3722 2904 -1698 2906
rect -1644 2904 -1631 2958
rect 22384 2948 28676 2992
rect 22384 2922 28326 2948
rect -1698 2894 -1644 2904
rect -5184 2824 -5178 2876
rect -5126 2871 -5120 2876
rect -4436 2871 -4430 2876
rect -5126 2829 -4430 2871
rect -5126 2824 -5120 2829
rect -4436 2824 -4430 2829
rect -4378 2824 -4372 2876
rect -3870 2798 -3864 2850
rect -3812 2848 -3806 2850
rect -1506 2848 -1500 2850
rect -3812 2800 -1500 2848
rect -3812 2798 -3806 2800
rect -1506 2798 -1500 2800
rect -1448 2798 -1442 2850
rect -871 2842 -862 2902
rect -802 2898 -793 2902
rect -802 2846 9928 2898
rect 9980 2846 9986 2898
rect -802 2842 -793 2846
rect -5416 2762 -5332 2776
rect -3670 2762 -3618 2768
rect -6006 2710 -6000 2762
rect -5948 2758 -5942 2762
rect -5416 2758 -5398 2762
rect -5948 2714 -5398 2758
rect -5948 2710 -5942 2714
rect -5416 2710 -5398 2714
rect -5346 2758 -5332 2762
rect -4804 2758 -4798 2762
rect -5346 2714 -4798 2758
rect -5346 2710 -5332 2714
rect -4804 2710 -4798 2714
rect -4746 2758 -4740 2762
rect -4746 2714 -3670 2758
rect -4746 2710 -4740 2714
rect 489 2731 495 2797
rect 561 2731 12415 2797
rect 12481 2731 12487 2797
rect 12988 2770 12994 2822
rect 13046 2770 13660 2822
rect 13712 2770 13718 2822
rect -5416 2692 -5332 2710
rect -3670 2704 -3618 2710
rect -3508 2614 -3502 2666
rect -3450 2657 -3444 2666
rect -2677 2657 -2671 2666
rect -3450 2623 -2671 2657
rect -3450 2614 -3444 2623
rect -2677 2614 -2671 2623
rect -2619 2614 -2613 2666
rect -1001 2645 -995 2703
rect -937 2645 11195 2703
rect 11253 2645 11259 2703
rect 13138 2631 13144 2686
rect 13199 2631 13788 2686
rect 13843 2631 13849 2686
rect 22384 2658 22442 2922
rect 22858 2666 28326 2922
rect 28650 2666 28676 2948
rect 22858 2658 28676 2666
rect 22384 2622 28676 2658
rect 7060 2553 12759 2564
rect 6281 2483 6287 2553
rect 6357 2494 12759 2553
rect 12829 2494 12881 2564
rect 6357 2483 7153 2494
rect -4042 2416 -4028 2480
rect -3964 2470 -2376 2480
rect -3964 2418 -2914 2470
rect -2862 2418 -2428 2470
rect -3964 2416 -2376 2418
rect -4042 2408 -2376 2416
rect 6828 2230 6886 2240
rect -4216 1880 -4210 1952
rect -4138 1942 -2534 1952
rect -4138 1890 -2756 1942
rect -2704 1890 -2586 1942
rect -1506 1894 -1500 1946
rect -1448 1944 -1442 1946
rect 4754 1944 4760 1946
rect -1448 1896 4760 1944
rect -1448 1894 -1442 1896
rect 4754 1894 4760 1896
rect 4812 1894 4818 1946
rect -4138 1880 -2534 1890
rect 1888 1754 1894 1826
rect 1966 1754 3450 1826
rect 3522 1754 3528 1826
rect -3191 1659 -3185 1717
rect -3127 1659 1525 1717
rect 1583 1659 1589 1717
rect 6828 1608 6886 1618
rect 7088 2230 7142 2483
rect 7088 1608 7142 1618
rect 7344 2230 7402 2240
rect 7344 1608 7402 1618
rect 7604 2230 7658 2240
rect -4436 1538 -4430 1590
rect -4378 1585 -4372 1590
rect -2530 1585 -2524 1590
rect -4378 1543 -2524 1585
rect -4378 1538 -4372 1543
rect -2530 1538 -2524 1543
rect -2472 1538 -2466 1590
rect 2630 1526 2636 1578
rect 2688 1577 2694 1578
rect 5512 1577 5518 1578
rect 2688 1527 5518 1577
rect 2688 1526 2694 1527
rect 5512 1526 5518 1527
rect 5570 1526 5576 1578
rect 7604 1471 7658 1618
rect 7860 2230 7918 2240
rect 7860 1608 7918 1618
rect 8120 2230 8174 2240
rect 8120 1471 8174 1618
rect 8376 2230 8434 2240
rect 8376 1608 8434 1618
rect 8636 2230 8690 2494
rect 8636 1608 8690 1618
rect 8892 2230 8950 2240
rect 8892 1608 8950 1618
rect 9152 2230 9206 2494
rect 9152 1608 9206 1618
rect 9408 2230 9466 2240
rect 9408 1608 9466 1618
rect 9668 2230 9722 2240
rect 9668 1471 9722 1618
rect 9924 2230 9982 2240
rect 9924 1608 9982 1618
rect 10184 2230 10238 2240
rect 10184 1471 10238 1618
rect 10440 2230 10498 2240
rect 10440 1608 10498 1618
rect 10700 2230 10754 2494
rect 10700 1608 10754 1618
rect 10956 2230 11014 2240
rect 10956 1608 11014 1618
rect 11216 2230 11270 2494
rect 11216 1608 11270 1618
rect 11472 2230 11530 2240
rect 11472 1608 11530 1618
rect 11732 2230 11786 2240
rect 11732 1471 11786 1618
rect 11988 2230 12046 2240
rect 11988 1608 12046 1618
rect 12248 2230 12302 2240
rect 12248 1471 12302 1618
rect 12504 2230 12562 2240
rect 12504 1608 12562 1618
rect 12764 2230 12818 2494
rect 13914 2416 13920 2468
rect 13972 2467 13978 2468
rect 14694 2467 14700 2468
rect 13972 2417 14700 2467
rect 13972 2416 13978 2417
rect 14694 2416 14700 2417
rect 14752 2416 14758 2468
rect 16570 2372 16576 2424
rect 16628 2423 16634 2424
rect 17684 2423 17690 2424
rect 16628 2373 17690 2423
rect 16628 2372 16634 2373
rect 17684 2372 17690 2373
rect 17742 2372 17748 2424
rect 17905 2355 17911 2421
rect 17977 2355 22555 2421
rect 22621 2355 22627 2421
rect 12764 1608 12818 1618
rect 13020 2230 13078 2240
rect 18624 2152 18748 2154
rect 14524 2147 18748 2152
rect 14524 2142 17911 2147
rect 14652 2090 14782 2142
rect 14910 2090 15040 2142
rect 15168 2090 15298 2142
rect 15426 2090 15556 2142
rect 15684 2090 15814 2142
rect 15942 2090 16588 2142
rect 16718 2090 16846 2142
rect 16976 2090 17102 2142
rect 17232 2090 17911 2142
rect 14524 2081 17911 2090
rect 17977 2144 18748 2147
rect 17977 2090 18624 2144
rect 17977 2081 18748 2090
rect 14524 2080 18748 2081
rect 30836 2032 30842 2092
rect 30902 2032 32006 2092
rect 32066 2032 32072 2092
rect 33947 2006 34033 2010
rect 32708 1910 32714 2006
rect 32810 2001 34038 2006
rect 32810 1915 33947 2001
rect 34033 1915 34038 2001
rect 32810 1910 34038 1915
rect 33947 1906 34033 1910
rect 32848 1654 32854 1750
rect 32950 1745 34298 1750
rect 32950 1659 34207 1745
rect 34293 1659 34302 1745
rect 32950 1654 34298 1659
rect 13020 1608 13078 1618
rect -5846 1457 -5794 1463
rect -5184 1452 -5178 1457
rect -5794 1410 -5178 1452
rect -5184 1405 -5178 1410
rect -5126 1405 -5120 1457
rect -4582 1448 -4530 1454
rect -5846 1399 -5794 1405
rect -3870 1446 -3864 1448
rect -4530 1398 -3864 1446
rect -3870 1396 -3864 1398
rect -3812 1396 -3806 1448
rect -4582 1390 -4530 1396
rect 2410 1380 2416 1436
rect 2472 1380 5378 1436
rect 5434 1380 5440 1436
rect 6035 1392 6041 1471
rect 6120 1392 12960 1471
rect 13300 1457 13352 1463
rect 13653 1454 13662 1461
rect 13352 1408 13662 1454
rect 13300 1399 13352 1405
rect 13653 1401 13662 1408
rect 13722 1401 13731 1461
rect 6828 1244 6886 1254
rect 4898 1186 5010 1196
rect 6080 1182 6376 1192
rect 5010 1079 6080 1181
rect 6080 1068 6376 1078
rect 4898 866 5010 876
rect -5889 670 -5831 676
rect -5831 612 -5137 670
rect -5079 612 -5073 670
rect -4621 660 -4563 666
rect -5889 606 -5831 612
rect -4563 602 -3185 660
rect -3127 602 -3121 660
rect 6828 622 6886 632
rect 7088 1242 7142 1392
rect 7088 620 7142 630
rect 7344 1244 7402 1254
rect 7344 622 7402 632
rect 7604 1244 7658 1254
rect -4621 596 -4563 602
rect 7604 352 7658 632
rect 7860 1244 7918 1254
rect 7860 622 7918 632
rect 8120 1244 8174 1254
rect 8120 352 8174 632
rect 8376 1244 8434 1254
rect 8376 622 8434 632
rect 8636 1244 8690 1392
rect 8636 622 8690 632
rect 8892 1244 8950 1254
rect 8892 622 8950 632
rect 9152 1244 9206 1392
rect 9152 622 9206 632
rect 9408 1244 9466 1254
rect 9408 622 9466 632
rect 9668 1244 9722 1254
rect 9668 352 9722 632
rect 9924 1246 9980 1256
rect 9924 620 9980 630
rect 10184 1244 10238 1254
rect 10184 352 10238 632
rect 10440 1244 10498 1254
rect 10440 622 10498 632
rect 10700 1244 10754 1392
rect 10700 622 10754 632
rect 10956 1244 11014 1254
rect 10956 622 11014 632
rect 11216 1244 11270 1392
rect 11216 622 11270 632
rect 11472 1244 11530 1254
rect 11472 622 11530 632
rect 11732 1244 11786 1254
rect 11732 352 11786 632
rect 11988 1244 12046 1254
rect 11988 622 12046 632
rect 12248 1244 12302 1254
rect 12248 352 12302 632
rect 12504 1244 12562 1254
rect 12504 622 12562 632
rect 12764 1244 12818 1392
rect 12764 622 12818 632
rect 13020 1244 13078 1254
rect 19467 1035 22419 1037
rect 16722 961 16728 1035
rect 16802 1012 19581 1035
rect 16802 961 17690 1012
rect 17684 960 17690 961
rect 17742 961 19581 1012
rect 19655 961 22419 1035
rect 17742 960 17748 961
rect 19467 951 22419 961
rect 22505 951 22511 1037
rect 15914 806 15920 878
rect 15992 806 21580 878
rect 21652 806 21658 878
rect 13914 638 13920 690
rect 13972 689 13978 690
rect 15160 689 15166 690
rect 13972 639 15166 689
rect 13972 638 13978 639
rect 15160 638 15166 639
rect 15218 638 15224 690
rect 13020 622 13078 632
rect 6281 282 6287 352
rect 6357 282 12510 352
rect 5326 114 5438 116
rect 5512 114 5518 166
rect 5570 165 5576 166
rect 7889 165 7895 166
rect 5570 115 7895 165
rect 5570 114 5576 115
rect 7889 114 7895 115
rect 7947 114 7953 166
rect 5266 106 5438 114
rect 5266 104 5326 106
rect 5438 64 6914 74
rect 5438 -2 5832 64
rect 10959 1 10965 103
rect 11067 98 13517 103
rect 11067 6 13420 98
rect 13512 6 13521 98
rect 11067 1 13517 6
rect 5438 -10 6914 -2
rect -4672 -108 -4618 -102
rect 5370 -12 6914 -10
rect 5370 -20 5438 -12
rect -5850 -128 -5798 -122
rect -5242 -134 -5236 -128
rect -5798 -174 -5236 -134
rect -5242 -180 -5236 -174
rect -5184 -180 -5178 -128
rect -4618 -162 -4267 -108
rect -4213 -162 -4207 -108
rect 5266 -118 5370 -108
rect -4672 -168 -4618 -162
rect -5850 -186 -5798 -180
rect 2864 -296 4748 -286
rect 2864 -348 2902 -296
rect 2958 -348 3072 -296
rect 3274 -348 3388 -296
rect 3590 -348 3704 -296
rect 3906 -348 4020 -296
rect 4076 -348 4748 -296
rect 2864 -358 4748 -348
rect 4820 -358 4826 -286
rect 30744 -340 30753 -331
rect 3100 -414 3152 -408
rect -3961 -521 -3955 -447
rect -3881 -521 -3241 -447
rect -3167 -521 -3161 -447
rect 1348 -448 1510 -438
rect 2862 -454 3100 -416
rect 1510 -464 3100 -454
rect 1510 -502 2910 -464
rect 3220 -466 3226 -414
rect 3882 -418 4918 -408
rect 3100 -472 3152 -466
rect 4004 -476 4918 -418
rect 3882 -484 4918 -476
rect 4994 -484 5000 -408
rect 22413 -426 22419 -340
rect 22505 -350 30753 -340
rect 30839 -340 30848 -331
rect 30839 -350 31120 -340
rect 22505 -416 22996 -350
rect 22505 -417 30753 -416
rect 30839 -417 31120 -416
rect 22505 -426 31120 -417
rect 33654 -472 33762 -464
rect 3882 -486 4004 -484
rect 1348 -512 1510 -502
rect -3740 -588 -3636 -578
rect 22022 -608 22028 -528
rect 22108 -608 28020 -528
rect 30739 -568 30748 -472
rect 30844 -477 33762 -472
rect 30844 -563 33665 -477
rect 33751 -563 33762 -477
rect 30844 -568 33762 -563
rect 33654 -574 33762 -568
rect -3740 -678 -3636 -668
rect 2250 -722 2256 -670
rect 2308 -671 2314 -670
rect 5088 -671 5094 -670
rect 2308 -721 5094 -671
rect 2308 -722 2314 -721
rect 5088 -722 5094 -721
rect 5146 -722 5152 -670
rect 21847 -756 21853 -677
rect 21932 -756 24920 -677
rect -4634 -792 -4582 -786
rect -4582 -844 -4132 -792
rect -4080 -844 -4074 -792
rect -4634 -850 -4582 -844
rect -5803 -874 -5717 -868
rect -5717 -960 -5365 -874
rect -5279 -960 -5273 -874
rect -3247 -876 -3241 -802
rect -3167 -812 3862 -802
rect -3167 -866 -2336 -812
rect -2092 -866 -1878 -812
rect -1634 -866 -504 -812
rect -260 -866 -46 -812
rect 198 -866 412 -812
rect 656 -866 870 -812
rect 1114 -866 1328 -812
rect 1572 -866 1786 -812
rect 2030 -866 2244 -812
rect 2488 -866 2702 -812
rect 2946 -866 3160 -812
rect 3404 -866 3618 -812
rect 13520 -830 13526 -758
rect 13598 -768 21112 -758
rect 13598 -820 14524 -768
rect 14648 -820 14782 -768
rect 14906 -820 15040 -768
rect 15164 -820 15298 -768
rect 15422 -820 15556 -768
rect 15680 -820 15814 -768
rect 15938 -820 16072 -768
rect 16196 -820 16330 -768
rect 16454 -820 16588 -768
rect 16712 -820 16846 -768
rect 16970 -820 17104 -768
rect 17228 -820 17362 -768
rect 17486 -820 18136 -768
rect 18260 -820 18394 -768
rect 18518 -820 18652 -768
rect 18776 -820 18910 -768
rect 19034 -820 19168 -768
rect 19292 -820 19426 -768
rect 19550 -820 19684 -768
rect 19808 -820 19942 -768
rect 20066 -820 20200 -768
rect 20324 -820 20458 -768
rect 20582 -820 20716 -768
rect 20840 -820 20974 -768
rect 21098 -820 21112 -768
rect 13598 -830 21112 -820
rect 24841 -824 24920 -756
rect -3167 -876 3862 -866
rect 21696 -896 21702 -824
rect 21774 -896 22852 -824
rect -5803 -966 -5717 -960
rect -4341 -1036 -4332 -960
rect -4256 -1036 -3584 -960
rect -3458 -970 -1956 -960
rect -3458 -1026 -2014 -970
rect -3458 -1036 -1956 -1026
rect -182 -970 2090 -960
rect -124 -1026 734 -970
rect 792 -1026 1650 -970
rect 1708 -1026 2090 -970
rect -182 -1036 2090 -1026
rect 2166 -970 3540 -960
rect 2166 -1026 2566 -970
rect 2624 -1026 3482 -970
rect 2166 -1036 3540 -1026
rect 4746 -1054 4822 -1044
rect 22780 -1048 22852 -896
rect 24840 -900 24920 -824
rect 27940 -900 28020 -608
rect 31037 -900 31108 -833
rect 23822 -910 25946 -900
rect 25936 -966 25946 -910
rect 23822 -976 25946 -966
rect 26918 -910 29032 -900
rect 26918 -976 29032 -966
rect 30014 -910 33326 -900
rect 32128 -966 33326 -910
rect 30014 -976 33326 -966
rect 33402 -976 33408 -900
rect -3738 -1132 -3644 -1122
rect -3738 -1218 -3644 -1208
rect 4822 -1064 13018 -1054
rect 4822 -1068 7468 -1064
rect 4822 -1120 5920 -1068
rect 6052 -1120 6178 -1068
rect 6310 -1070 7468 -1068
rect 6310 -1120 6436 -1070
rect 4822 -1122 6436 -1120
rect 6568 -1074 7468 -1070
rect 6568 -1122 6694 -1074
rect 4822 -1130 6694 -1122
rect 6826 -1120 7468 -1074
rect 7600 -1120 7726 -1064
rect 7858 -1120 7984 -1064
rect 8116 -1120 8242 -1064
rect 8374 -1120 9016 -1064
rect 9148 -1120 9274 -1064
rect 9406 -1120 9532 -1064
rect 9664 -1120 9790 -1064
rect 9922 -1120 10048 -1064
rect 10180 -1120 10306 -1064
rect 10438 -1120 10564 -1064
rect 10696 -1120 10822 -1064
rect 10954 -1120 11080 -1064
rect 11212 -1120 11338 -1064
rect 11470 -1120 11596 -1064
rect 11728 -1120 11854 -1064
rect 11986 -1120 12112 -1064
rect 12244 -1120 12370 -1064
rect 12502 -1120 12628 -1064
rect 12760 -1120 12886 -1064
rect 22624 -1058 32294 -1048
rect 22748 -1110 22882 -1058
rect 23006 -1110 23656 -1058
rect 23780 -1110 23914 -1058
rect 24038 -1110 24172 -1058
rect 24296 -1110 24430 -1058
rect 24554 -1110 24688 -1058
rect 24812 -1110 24946 -1058
rect 25070 -1110 25204 -1058
rect 25328 -1110 25462 -1058
rect 25586 -1110 25718 -1058
rect 25842 -1110 25978 -1058
rect 26102 -1110 26752 -1058
rect 26876 -1110 27008 -1058
rect 27132 -1110 27268 -1058
rect 27392 -1110 27526 -1058
rect 27650 -1110 27784 -1058
rect 27908 -1110 28042 -1058
rect 28166 -1110 28300 -1058
rect 28424 -1110 28558 -1058
rect 28682 -1110 28816 -1058
rect 28940 -1110 29074 -1058
rect 29198 -1110 29848 -1058
rect 29972 -1110 30106 -1058
rect 30230 -1110 30364 -1058
rect 30488 -1110 30622 -1058
rect 30746 -1110 30880 -1058
rect 31004 -1110 31138 -1058
rect 31262 -1110 31396 -1058
rect 31520 -1110 31654 -1058
rect 31778 -1110 31912 -1058
rect 32036 -1110 32170 -1058
rect 22624 -1120 32294 -1110
rect 6826 -1130 13018 -1120
rect 6436 -1132 6568 -1130
rect 6694 -1140 6826 -1130
rect 19518 -1208 19698 -1198
rect 14688 -1218 19518 -1208
rect 13976 -1224 13982 -1218
rect 4950 -1282 5027 -1276
rect 13782 -1279 13788 -1224
rect 13843 -1270 13982 -1224
rect 14034 -1224 14040 -1218
rect 14034 -1270 14688 -1224
rect 14742 -1270 16236 -1218
rect 16290 -1270 16752 -1218
rect 16806 -1270 18300 -1218
rect 18354 -1270 18816 -1218
rect 18870 -1270 19518 -1218
rect 13843 -1279 19518 -1270
rect 14688 -1280 19518 -1279
rect 19698 -1218 20418 -1208
rect 19698 -1270 20364 -1218
rect 19698 -1280 20418 -1270
rect 4822 -1300 4950 -1282
rect 4746 -1310 4950 -1300
rect 4748 -1358 4950 -1310
rect 4748 -1525 4820 -1358
rect 5027 -1286 13601 -1282
rect 5027 -1357 13527 -1286
rect 13598 -1357 13604 -1286
rect 19518 -1290 19698 -1280
rect 5027 -1359 13601 -1357
rect 4950 -1365 5027 -1359
rect 15924 -1374 16076 -1368
rect 15204 -1378 19900 -1374
rect 15204 -1384 15924 -1378
rect 13654 -1438 13660 -1386
rect 13712 -1436 15204 -1386
rect 15258 -1436 15720 -1384
rect 15774 -1436 15924 -1384
rect 13712 -1438 15924 -1436
rect 15204 -1446 15924 -1438
rect 16076 -1384 19900 -1378
rect 16076 -1436 17268 -1384
rect 17322 -1436 17784 -1384
rect 17838 -1436 19332 -1384
rect 19386 -1436 19846 -1384
rect 16076 -1446 19900 -1436
rect 15924 -1460 16076 -1450
rect 4726 -1602 4732 -1525
rect 4809 -1602 4950 -1525
rect 5027 -1602 5033 -1525
rect 6808 -1608 7774 -1602
rect 6808 -1614 13096 -1608
rect -4691 -1687 -4685 -1625
rect -4623 -1687 -3235 -1625
rect -3173 -1687 -3167 -1625
rect 6202 -1674 6208 -1622
rect 6260 -1625 6266 -1622
rect 6808 -1625 6824 -1614
rect 6260 -1671 6824 -1625
rect 6260 -1674 6266 -1671
rect 6808 -1686 6824 -1671
rect 6890 -1686 7340 -1614
rect 7406 -1686 7856 -1614
rect 7922 -1686 8888 -1614
rect 8954 -1686 9920 -1614
rect 9986 -1686 10952 -1614
rect 11018 -1618 11984 -1614
rect 11018 -1686 11680 -1618
rect 11882 -1686 11984 -1618
rect 12050 -1686 12500 -1614
rect 12566 -1686 13016 -1614
rect 13082 -1686 13096 -1614
rect 6808 -1694 13096 -1686
rect 11680 -1696 11882 -1694
rect -5888 -1704 -5822 -1700
rect -5486 -1704 -5410 -1696
rect -5888 -1709 -5479 -1704
rect -5888 -1761 -5880 -1709
rect -5828 -1761 -5479 -1709
rect -5888 -1766 -5479 -1761
rect -5417 -1766 -5410 -1704
rect -5888 -1768 -5822 -1766
rect -5486 -1774 -5410 -1766
rect 8148 -1728 8406 -1724
rect 11474 -1728 11528 -1724
rect 8148 -1734 11528 -1728
rect 8406 -1738 11474 -1734
rect 8432 -1786 11474 -1738
rect 8432 -1790 11528 -1786
rect 8406 -1796 11528 -1790
rect 22534 -1796 22600 -1786
rect 8406 -1800 8432 -1796
rect 8148 -1810 8406 -1800
rect -3284 -1834 -3204 -1824
rect -3204 -1844 -1496 -1834
rect 22528 -1838 22534 -1798
rect -3204 -1904 -2474 -1844
rect -2412 -1904 -1558 -1844
rect 23050 -1796 23116 -1786
rect 22600 -1838 23050 -1798
rect 22534 -1878 22600 -1868
rect 25630 -1792 25696 -1782
rect 31040 -1786 31104 -1776
rect 23116 -1838 25630 -1798
rect 28728 -1796 28792 -1786
rect 25696 -1838 28728 -1798
rect 23050 -1878 23116 -1868
rect 24588 -1878 24674 -1868
rect -3204 -1914 -1496 -1904
rect 21862 -1894 21932 -1882
rect -3284 -1926 -3204 -1916
rect 21862 -1946 21871 -1894
rect 21923 -1908 21932 -1894
rect 24588 -1908 24598 -1878
rect 21923 -1946 24598 -1908
rect 21862 -1950 24598 -1946
rect 24664 -1899 24674 -1878
rect 25114 -1878 25180 -1868
rect 25630 -1874 25696 -1864
rect 28792 -1838 31040 -1798
rect 31308 -1792 31368 -1782
rect 31104 -1838 31308 -1798
rect 31040 -1858 31104 -1848
rect 31824 -1792 31884 -1782
rect 31368 -1838 31824 -1798
rect 28728 -1868 28792 -1858
rect 31308 -1864 31368 -1854
rect 31884 -1838 32184 -1798
rect 31824 -1864 31884 -1854
rect 24664 -1906 24856 -1899
rect 24664 -1946 25114 -1906
rect 24664 -1950 24674 -1946
rect 21862 -1952 24674 -1950
rect 21862 -1958 21932 -1952
rect -4422 -2023 -4416 -1958
rect -4351 -2023 -3100 -1958
rect -3035 -2023 -3029 -1958
rect 24588 -1960 24674 -1952
rect 26146 -1878 26212 -1868
rect 25180 -1946 26146 -1906
rect 25114 -1960 25180 -1950
rect 27942 -1898 28010 -1888
rect 26212 -1946 27942 -1906
rect 26146 -1960 26212 -1950
rect 28210 -1902 28274 -1892
rect 28010 -1946 28210 -1906
rect 27942 -1964 28010 -1954
rect 29244 -1900 29304 -1890
rect 28274 -1946 29244 -1906
rect 28210 -1974 28274 -1964
rect 29760 -1898 29820 -1888
rect 29304 -1946 29760 -1906
rect 29244 -1972 29304 -1962
rect 29820 -1946 29832 -1906
rect 29760 -1970 29820 -1960
rect 23566 -1992 23632 -1982
rect 23562 -2048 23566 -2004
rect 24082 -1992 24148 -1982
rect 23632 -2048 24082 -2004
rect 23566 -2074 23632 -2064
rect 24850 -2000 24908 -1990
rect 24148 -2048 24850 -2004
rect 26662 -1992 26728 -1982
rect 24908 -2048 26662 -2004
rect 24850 -2062 24908 -2052
rect 24082 -2074 24148 -2064
rect 26728 -2018 30880 -2004
rect 26728 -2020 30274 -2018
rect 26728 -2048 27696 -2020
rect 26662 -2074 26728 -2064
rect 27760 -2048 30274 -2020
rect 27174 -2094 27250 -2084
rect 27696 -2092 27760 -2082
rect 30338 -2048 30792 -2018
rect 30274 -2090 30338 -2080
rect 30856 -2048 30880 -2018
rect 30792 -2090 30856 -2080
rect -2474 -2166 -2412 -2162
rect -1558 -2166 -1496 -2160
rect -642 -2166 -580 -2160
rect 256 -2166 352 -2164
rect 1190 -2166 1252 -2160
rect 3942 -2164 4022 -2154
rect -3113 -2244 -3107 -2166
rect -3029 -2170 3942 -2166
rect -3029 -2172 -1558 -2170
rect -3029 -2234 -2474 -2172
rect -2412 -2232 -1558 -2172
rect -1496 -2232 -642 -2170
rect -580 -2174 1190 -2170
rect -580 -2232 256 -2174
rect -2412 -2234 256 -2232
rect -3029 -2242 256 -2234
rect 352 -2232 1190 -2174
rect 1252 -2176 3942 -2170
rect 1252 -2232 2106 -2176
rect 352 -2238 2106 -2232
rect 2168 -2178 3942 -2176
rect 2168 -2232 3026 -2178
rect 3080 -2232 3942 -2178
rect 2168 -2238 3942 -2232
rect 352 -2242 3942 -2238
rect -3029 -2244 3942 -2242
rect 27174 -2174 27250 -2164
rect 256 -2252 352 -2244
rect 2106 -2248 2168 -2244
rect 3942 -2254 4022 -2244
rect -3736 -2264 -3640 -2254
rect -3736 -2366 -3640 -2356
rect -5886 -2481 -5816 -2472
rect -5886 -2533 -5875 -2481
rect -5823 -2486 -5816 -2481
rect -5590 -2486 -5584 -2481
rect -5823 -2528 -5584 -2486
rect -5823 -2533 -5816 -2528
rect -5590 -2533 -5584 -2528
rect -5532 -2533 -5526 -2481
rect -5886 -2542 -5816 -2533
rect 4688 -2614 4798 -2604
rect 5088 -2627 5094 -2626
rect 4798 -2677 5094 -2627
rect 5088 -2678 5094 -2677
rect 5146 -2678 5152 -2626
rect 4688 -2700 4798 -2690
rect -3738 -2818 -3642 -2808
rect 21580 -2910 21652 -2904
rect -3738 -2920 -3642 -2910
rect 14524 -2920 21580 -2910
rect 260 -2962 348 -2952
rect -3282 -3038 -3202 -3028
rect 258 -3042 260 -2974
rect -3202 -3108 260 -3042
rect 20582 -2972 21580 -2920
rect 348 -3108 354 -2974
rect 14524 -2982 21580 -2972
rect 21580 -2988 21652 -2982
rect 22634 -2952 31798 -2942
rect 22758 -2953 22892 -2952
rect 22758 -3006 22817 -2953
rect 22634 -3011 22817 -3006
rect 22875 -3006 22892 -2953
rect 23016 -3006 23150 -2952
rect 23274 -3006 23408 -2952
rect 23532 -3006 23666 -2952
rect 23790 -3006 23924 -2952
rect 24048 -3006 24696 -2952
rect 24820 -3006 24956 -2952
rect 25080 -3006 25216 -2952
rect 25340 -3006 25474 -2952
rect 25598 -3006 25730 -2952
rect 25854 -3006 25988 -2952
rect 26112 -2954 30374 -2952
rect 26112 -3006 26244 -2954
rect 22875 -3008 26244 -3006
rect 26368 -3008 26506 -2954
rect 26630 -3008 26762 -2954
rect 26886 -3008 27022 -2954
rect 27404 -3008 27538 -2954
rect 27662 -3008 27794 -2954
rect 27918 -2956 28310 -2954
rect 27918 -3008 28054 -2956
rect 22875 -3010 28054 -3008
rect 28178 -3008 28310 -2956
rect 28434 -3008 28568 -2954
rect 28692 -3008 28826 -2954
rect 28950 -3008 29084 -2954
rect 29208 -3008 29342 -2954
rect 29466 -3008 29600 -2954
rect 29724 -3006 30374 -2954
rect 30498 -3006 30632 -2952
rect 30756 -3006 30890 -2952
rect 31014 -3006 31148 -2952
rect 31272 -3006 31406 -2952
rect 31530 -3006 31664 -2952
rect 31788 -3006 31798 -2952
rect 29724 -3008 31798 -3006
rect 28178 -3010 31798 -3008
rect 22875 -3011 31798 -3010
rect 22634 -3016 31798 -3011
rect 26244 -3018 26368 -3016
rect 26506 -3018 26630 -3016
rect 26762 -3018 26886 -3016
rect 27022 -3018 27404 -3016
rect 27538 -3018 27662 -3016
rect 27794 -3018 27918 -3016
rect 28054 -3020 28178 -3016
rect 28310 -3018 28434 -3016
rect 28568 -3018 28692 -3016
rect 28826 -3018 28950 -3016
rect 29084 -3018 29208 -3016
rect 29342 -3018 29466 -3016
rect 29600 -3018 29724 -3016
rect -3202 -3112 354 -3108
rect 5290 -3040 5482 -3030
rect -3202 -3114 352 -3112
rect 260 -3118 348 -3114
rect -3282 -3130 -3202 -3120
rect 10532 -3054 10664 -3050
rect 5482 -3064 12986 -3054
rect 5482 -3124 6920 -3064
rect 9364 -3124 9510 -3064
rect 10396 -3124 10546 -3064
rect 5482 -3134 12986 -3124
rect 10184 -3136 10408 -3134
rect 5290 -3156 5482 -3146
rect 6326 -3180 6388 -3178
rect 9410 -3180 9464 -3178
rect 10442 -3180 10496 -3178
rect -886 -3190 -792 -3184
rect 6313 -3188 10496 -3180
rect -5876 -3285 -5824 -3279
rect -5696 -3288 -5690 -3285
rect -5824 -3334 -5690 -3288
rect -5696 -3337 -5690 -3334
rect -5638 -3337 -5632 -3285
rect -4697 -3300 -4691 -3190
rect -4581 -3300 -3955 -3190
rect -3845 -3194 2868 -3190
rect -3845 -3202 -886 -3194
rect -3845 -3204 -1340 -3202
rect -3845 -3290 -2264 -3204
rect -2170 -3290 -1804 -3204
rect -1710 -3288 -1340 -3204
rect -1246 -3280 -886 -3202
rect -792 -3202 2868 -3194
rect -792 -3204 1398 -3202
rect -792 -3280 -432 -3204
rect -1246 -3288 -432 -3280
rect -1710 -3290 -432 -3288
rect -338 -3290 30 -3204
rect 124 -3206 948 -3204
rect 124 -3290 482 -3206
rect -3845 -3292 482 -3290
rect 576 -3290 948 -3206
rect 1042 -3288 1398 -3204
rect 1492 -3204 2314 -3202
rect 1492 -3288 1856 -3204
rect 1042 -3290 1856 -3288
rect 1950 -3288 2314 -3204
rect 2408 -3204 2868 -3202
rect 2408 -3288 2770 -3204
rect 1950 -3290 2770 -3288
rect 2864 -3290 2868 -3204
rect 6313 -3242 6326 -3188
rect 6388 -3240 9410 -3188
rect 9464 -3240 10442 -3188
rect 6388 -3242 10496 -3240
rect 9410 -3250 9464 -3242
rect 10442 -3250 10496 -3242
rect 6326 -3260 6388 -3250
rect 576 -3292 2868 -3290
rect -3845 -3298 2868 -3292
rect -3845 -3300 -2170 -3298
rect -1804 -3300 -1710 -3298
rect -432 -3300 -338 -3298
rect 30 -3300 124 -3298
rect 482 -3302 576 -3298
rect 948 -3300 1042 -3298
rect 1856 -3300 1950 -3298
rect 2770 -3300 2864 -3298
rect -5876 -3343 -5824 -3337
rect -4138 -3510 -4132 -3458
rect -4080 -3510 5320 -3458
rect 5372 -3510 5378 -3458
rect -4267 -3543 14682 -3542
rect -4273 -3597 -4267 -3543
rect -4213 -3597 14682 -3543
rect 14737 -3597 14743 -3542
rect -5480 -3762 -5474 -3710
rect -5422 -3713 -5416 -3710
rect 13656 -3713 13662 -3710
rect -5422 -3759 13662 -3713
rect -5422 -3762 -5416 -3759
rect 13656 -3762 13662 -3759
rect 13714 -3762 13720 -3710
rect -5590 -3876 -5584 -3824
rect -5532 -3829 -5526 -3824
rect 13976 -3829 13982 -3824
rect -5532 -3871 13982 -3829
rect -5532 -3876 -5526 -3871
rect 13976 -3876 13982 -3871
rect 14034 -3876 14040 -3824
rect -5690 -3920 -5638 -3914
rect 6202 -3923 6208 -3920
rect -5638 -3969 6208 -3923
rect 6202 -3972 6208 -3969
rect 6260 -3972 6266 -3920
rect -5690 -3978 -5638 -3972
rect -5364 -4102 -5358 -4029
rect -5285 -4102 21705 -4029
rect 21778 -4102 21784 -4029
rect -5242 -4268 -5236 -4216
rect -5184 -4223 -5178 -4216
rect 21864 -4221 21870 -4215
rect 1262 -4223 21870 -4221
rect -5184 -4261 21870 -4223
rect -5184 -4268 -5178 -4261
rect 1262 -4262 21870 -4261
rect 21864 -4267 21870 -4262
rect 21922 -4267 21928 -4215
rect -5143 -4399 -5137 -4341
rect -5079 -4399 22817 -4341
rect 22875 -4399 22881 -4341
<< via2 >>
rect -5190 13702 -5106 13786
rect 12478 12942 12550 13014
rect 13351 12951 13413 13013
rect 13346 12729 13418 12801
rect 22385 12153 22467 12235
rect 11330 11762 11418 11850
rect 13385 11797 13447 11859
rect 12483 11331 12545 11393
rect 13380 11328 13452 11400
rect 2702 10252 2758 10308
rect 2511 9482 2567 9538
rect 30582 8874 30678 8970
rect 33431 8879 33517 8965
rect 30587 8707 30673 8793
rect 2699 8479 2761 8541
rect 22380 7868 22472 7960
rect 9915 7393 10021 7499
rect -3775 7103 -3709 7169
rect 2336 7150 2392 7206
rect 2509 7007 2570 7068
rect 2836 6996 2892 7052
rect 2526 6828 2582 6884
rect 2834 6826 2894 6886
rect -3328 6236 -3272 6292
rect -4114 5494 -4058 5550
rect 3254 5394 3310 6616
rect 3770 5394 3826 6616
rect 4286 5394 4342 6616
rect 4802 5394 4858 6616
rect 5318 5394 5374 6616
rect 5834 5394 5890 6616
rect 6350 5394 6406 6616
rect 6866 5394 6922 6616
rect 7382 5394 7438 6616
rect 7898 5394 7954 6616
rect 8414 5394 8470 6616
rect 8930 5394 8986 6616
rect 9446 5394 9502 6616
rect -4327 4585 -4261 4651
rect -3780 4580 -3704 4656
rect 2524 4610 2584 4670
rect 3254 3790 3310 5012
rect 3770 3790 3826 5012
rect 4286 3790 4342 5012
rect 4802 3790 4858 5012
rect 5318 3790 5374 5012
rect 5834 3790 5890 5012
rect 6350 3790 6406 5012
rect 6866 3790 6922 5012
rect 7382 3790 7438 5012
rect 7898 3790 7954 5012
rect 8414 3790 8470 5012
rect 8930 3790 8986 5012
rect 9446 3790 9502 5012
rect 2332 3458 2396 3522
rect -4116 3000 -4056 3060
rect 13664 3002 13720 3058
rect -3720 2906 -3664 2962
rect -862 2842 -802 2902
rect 22442 2658 22858 2922
rect 6828 1618 6830 2230
rect 6830 1618 6884 2230
rect 6884 1618 6886 2230
rect 7344 1618 7346 2230
rect 7346 1618 7400 2230
rect 7400 1618 7402 2230
rect 7860 1618 7862 2230
rect 7862 1618 7916 2230
rect 7916 1618 7918 2230
rect 8376 1618 8378 2230
rect 8378 1618 8432 2230
rect 8432 1618 8434 2230
rect 8892 1618 8894 2230
rect 8894 1618 8948 2230
rect 8948 1618 8950 2230
rect 9408 1618 9410 2230
rect 9410 1618 9464 2230
rect 9464 1618 9466 2230
rect 9924 1618 9926 2230
rect 9926 1618 9980 2230
rect 9980 1618 9982 2230
rect 10440 1618 10442 2230
rect 10442 1618 10496 2230
rect 10496 1618 10498 2230
rect 10956 1618 10958 2230
rect 10958 1618 11012 2230
rect 11012 1618 11014 2230
rect 11472 1618 11474 2230
rect 11474 1618 11528 2230
rect 11528 1618 11530 2230
rect 11988 1618 11990 2230
rect 11990 1618 12044 2230
rect 12044 1618 12046 2230
rect 12504 1618 12506 2230
rect 12506 1618 12560 2230
rect 12560 1618 12562 2230
rect 13020 1618 13022 2230
rect 13022 1618 13076 2230
rect 13076 1618 13078 2230
rect 33947 1915 34033 2001
rect 34207 1659 34293 1745
rect 13662 1401 13722 1461
rect 6080 1078 6376 1182
rect 6828 632 6830 1244
rect 6830 632 6884 1244
rect 6884 632 6886 1244
rect 7344 632 7346 1244
rect 7346 632 7400 1244
rect 7400 632 7402 1244
rect 7860 632 7862 1244
rect 7862 632 7916 1244
rect 7916 632 7918 1244
rect 8376 632 8378 1244
rect 8378 632 8432 1244
rect 8432 632 8434 1244
rect 8892 632 8894 1244
rect 8894 632 8948 1244
rect 8948 632 8950 1244
rect 9408 632 9410 1244
rect 9410 632 9464 1244
rect 9464 632 9466 1244
rect 9924 632 9926 1246
rect 9926 632 9978 1246
rect 9978 632 9980 1246
rect 9924 630 9980 632
rect 10440 632 10442 1244
rect 10442 632 10496 1244
rect 10496 632 10498 1244
rect 10956 632 10958 1244
rect 10958 632 11012 1244
rect 11012 632 11014 1244
rect 11472 632 11474 1244
rect 11474 632 11528 1244
rect 11528 632 11530 1244
rect 11988 632 11990 1244
rect 11990 632 12044 1244
rect 12044 632 12046 1244
rect 12504 632 12506 1244
rect 12506 632 12560 1244
rect 12560 632 12562 1244
rect 13020 632 13022 1244
rect 13022 632 13076 1244
rect 13076 632 13078 1244
rect 13420 6 13512 98
rect 30753 -350 30839 -331
rect 30753 -416 30839 -350
rect 30753 -417 30839 -416
rect -3740 -668 -3636 -588
rect 30748 -568 30844 -472
rect 33665 -563 33751 -477
rect -4332 -1036 -4256 -960
rect -3738 -1208 -3644 -1132
rect -3736 -2356 -3640 -2264
rect -3738 -2910 -3642 -2818
<< metal3 >>
rect -5195 13786 -5101 13791
rect -5195 13702 -5190 13786
rect -5106 13784 -5101 13786
rect 11330 13784 11418 13788
rect -5106 13704 11422 13784
rect -5106 13702 -5101 13704
rect -5195 13697 -5101 13702
rect 11330 11855 11418 13704
rect 12473 13014 12555 13019
rect 12473 12942 12478 13014
rect 12550 12942 12555 13014
rect 12473 12937 12555 12942
rect 13346 13013 13418 13018
rect 13346 12951 13351 13013
rect 13413 12951 13418 13013
rect 11325 11850 11423 11855
rect 11325 11762 11330 11850
rect 11418 11762 11423 11850
rect 11325 11757 11423 11762
rect 12478 11393 12550 12937
rect 13346 12806 13418 12951
rect 13341 12801 13423 12806
rect 13341 12729 13346 12801
rect 13418 12729 13423 12801
rect 13341 12724 13423 12729
rect 33426 12499 33522 12542
rect 33423 12493 33525 12499
rect 33423 12385 33525 12391
rect 22380 12235 22472 12240
rect 22380 12153 22385 12235
rect 22467 12153 22472 12235
rect 13380 11859 13452 11864
rect 13380 11797 13385 11859
rect 13447 11797 13452 11859
rect 13380 11405 13452 11797
rect 12478 11331 12483 11393
rect 12545 11331 12550 11393
rect 12478 11326 12550 11331
rect 13375 11400 13457 11405
rect 13375 11328 13380 11400
rect 13452 11328 13457 11400
rect 13375 11323 13457 11328
rect 2697 10308 2763 10313
rect 2697 10252 2702 10308
rect 2758 10252 2763 10308
rect 2697 10247 2763 10252
rect 2506 9538 2572 9543
rect 2506 9482 2511 9538
rect 2567 9482 2572 9538
rect 2506 9477 2572 9482
rect 2331 7206 2397 7211
rect -3780 7169 -3704 7174
rect -3780 7103 -3775 7169
rect -3709 7103 -3704 7169
rect 2331 7150 2336 7206
rect 2392 7150 2397 7206
rect 2331 7145 2397 7150
rect -4119 5550 -4053 5555
rect -4119 5494 -4114 5550
rect -4058 5494 -4053 5550
rect -4119 5489 -4053 5494
rect -4332 4651 -4256 4656
rect -4332 4585 -4327 4651
rect -4261 4585 -4256 4651
rect -4332 -955 -4256 4585
rect -4116 3065 -4056 5489
rect -3780 4661 -3704 7103
rect -3333 6294 -3267 6297
rect -3333 6292 -802 6294
rect -3333 6236 -3328 6292
rect -3272 6236 -802 6292
rect -3333 6234 -802 6236
rect -3333 6231 -3267 6234
rect -3785 4656 -3699 4661
rect -3785 4580 -3780 4656
rect -3704 4580 -3699 4656
rect -3785 4575 -3699 4580
rect -4121 3060 -4051 3065
rect -4121 3000 -4116 3060
rect -4056 3000 -4051 3060
rect -4121 2995 -4051 3000
rect -3725 2962 -3659 2967
rect -3725 2906 -3720 2962
rect -3664 2906 -3659 2962
rect -862 2907 -802 6234
rect 2332 3527 2396 7145
rect 2508 7073 2570 9477
rect 2699 8546 2761 10247
rect 2694 8541 2766 8546
rect 2694 8479 2699 8541
rect 2761 8479 2766 8541
rect 2694 8474 2766 8479
rect 22380 7965 22472 12153
rect 30577 8970 30683 8975
rect 30577 8874 30582 8970
rect 30678 8874 30683 8970
rect 30577 8869 30683 8874
rect 33426 8965 33522 12385
rect 33660 9487 33756 12560
rect 33942 11019 34038 12542
rect 33941 11013 34043 11019
rect 33941 10905 34043 10911
rect 33653 9481 33756 9487
rect 33755 9379 33756 9481
rect 33653 9373 33756 9379
rect 33426 8879 33431 8965
rect 33517 8879 33522 8965
rect 30582 8793 30678 8869
rect 30582 8707 30587 8793
rect 30673 8707 30678 8793
rect 30582 8702 30678 8707
rect 22375 7960 22477 7965
rect 22375 7868 22380 7960
rect 22472 7868 22477 7960
rect 22375 7863 22477 7868
rect 9910 7499 10026 7504
rect 9910 7393 9915 7499
rect 10021 7393 10026 7499
rect 2504 7068 2575 7073
rect 2504 7007 2509 7068
rect 2570 7007 2575 7068
rect 2504 7002 2575 7007
rect 2831 7052 2897 7057
rect 2831 6996 2836 7052
rect 2892 6996 2897 7052
rect 2831 6991 2897 6996
rect 2834 6891 2894 6991
rect 2521 6884 2587 6889
rect 2521 6828 2526 6884
rect 2582 6828 2587 6884
rect 2521 6823 2587 6828
rect 2829 6886 2899 6891
rect 2829 6826 2834 6886
rect 2894 6826 2899 6886
rect 2524 4675 2584 6823
rect 2829 6821 2899 6826
rect 3244 6616 3320 6708
rect 3244 5394 3254 6616
rect 3310 5394 3320 6616
rect 3244 5264 3320 5394
rect 3760 6616 3836 6708
rect 3760 5394 3770 6616
rect 3826 5394 3836 6616
rect 3760 5264 3836 5394
rect 4276 6616 4352 6708
rect 4276 5394 4286 6616
rect 4342 5394 4352 6616
rect 4276 5264 4352 5394
rect 4792 6616 4868 6708
rect 4792 5394 4802 6616
rect 4858 5394 4868 6616
rect 4792 5264 4868 5394
rect 5308 6616 5384 6708
rect 5308 5394 5318 6616
rect 5374 5394 5384 6616
rect 5308 5264 5384 5394
rect 5824 6616 5900 6708
rect 5824 5394 5834 6616
rect 5890 5394 5900 6616
rect 5824 5264 5900 5394
rect 6340 6616 6416 6708
rect 6340 5394 6350 6616
rect 6406 5394 6416 6616
rect 6340 5264 6416 5394
rect 6856 6616 6932 6708
rect 6856 5394 6866 6616
rect 6922 5394 6932 6616
rect 6856 5264 6932 5394
rect 7372 6616 7448 6708
rect 7372 5394 7382 6616
rect 7438 5394 7448 6616
rect 7372 5264 7448 5394
rect 7888 6616 7964 6708
rect 7888 5394 7898 6616
rect 7954 5394 7964 6616
rect 7888 5264 7964 5394
rect 8404 6616 8480 6708
rect 8404 5394 8414 6616
rect 8470 5394 8480 6616
rect 8404 5264 8480 5394
rect 8920 6616 8996 6708
rect 8920 5394 8930 6616
rect 8986 5394 8996 6616
rect 8920 5264 8996 5394
rect 9436 6616 9512 6708
rect 9436 5394 9446 6616
rect 9502 5394 9512 6616
rect 9436 5264 9512 5394
rect 9910 5264 10026 7393
rect 33426 6475 33522 8879
rect 33417 6469 33522 6475
rect 33519 6367 33522 6469
rect 33417 6361 33522 6367
rect 3224 5148 10026 5264
rect 3244 5012 3320 5148
rect 2519 4670 2589 4675
rect 2519 4610 2524 4670
rect 2584 4610 2589 4670
rect 2519 4605 2589 4610
rect 3244 3790 3254 5012
rect 3310 3790 3320 5012
rect 3244 3770 3320 3790
rect 3760 5012 3836 5148
rect 3760 3790 3770 5012
rect 3826 3790 3836 5012
rect 3760 3770 3836 3790
rect 4276 5012 4352 5148
rect 4276 3790 4286 5012
rect 4342 3790 4352 5012
rect 4276 3770 4352 3790
rect 4792 5012 4868 5148
rect 4792 3790 4802 5012
rect 4858 3790 4868 5012
rect 4792 3770 4868 3790
rect 5308 5012 5384 5148
rect 5308 3790 5318 5012
rect 5374 3790 5384 5012
rect 5308 3770 5384 3790
rect 5824 5012 5900 5148
rect 5824 3790 5834 5012
rect 5890 3790 5900 5012
rect 5824 3770 5900 3790
rect 6340 5012 6416 5148
rect 6340 3790 6350 5012
rect 6406 3790 6416 5012
rect 6340 3770 6416 3790
rect 6856 5012 6932 5148
rect 6856 3790 6866 5012
rect 6922 3790 6932 5012
rect 6856 3770 6932 3790
rect 7372 5012 7448 5148
rect 7372 3790 7382 5012
rect 7438 3790 7448 5012
rect 7372 3770 7448 3790
rect 7888 5012 7964 5148
rect 7888 3790 7898 5012
rect 7954 3790 7964 5012
rect 7888 3770 7964 3790
rect 8404 5012 8480 5148
rect 8404 3790 8414 5012
rect 8470 3790 8480 5012
rect 8404 3770 8480 3790
rect 8920 5012 8996 5148
rect 8920 3790 8930 5012
rect 8986 3790 8996 5012
rect 8920 3770 8996 3790
rect 9436 5012 9512 5148
rect 9436 3790 9446 5012
rect 9502 3790 9512 5012
rect 9436 3770 9512 3790
rect 2327 3522 2401 3527
rect 2327 3458 2332 3522
rect 2396 3458 2401 3522
rect 2327 3453 2401 3458
rect 13659 3058 13725 3063
rect 13659 3002 13664 3058
rect 13720 3002 13725 3058
rect 13659 2997 13725 3002
rect -3725 2901 -3659 2906
rect -867 2902 -797 2907
rect -3722 -583 -3662 2901
rect -867 2842 -862 2902
rect -802 2842 -797 2902
rect -867 2837 -797 2842
rect 6818 2230 6896 2235
rect 6818 1618 6828 2230
rect 6886 1618 6896 2230
rect 6818 1482 6896 1618
rect 7334 2230 7412 2235
rect 7334 1618 7344 2230
rect 7402 1618 7412 2230
rect 7334 1482 7412 1618
rect 7850 2230 7928 2235
rect 7850 1618 7860 2230
rect 7918 1618 7928 2230
rect 7850 1482 7928 1618
rect 8366 2230 8444 2235
rect 8366 1618 8376 2230
rect 8434 1618 8444 2230
rect 8366 1482 8444 1618
rect 8882 2230 8960 2235
rect 8882 1618 8892 2230
rect 8950 1618 8960 2230
rect 8882 1482 8960 1618
rect 9398 2230 9476 2235
rect 9398 1618 9408 2230
rect 9466 1618 9476 2230
rect 9398 1482 9476 1618
rect 9914 2230 9992 2235
rect 9914 1618 9924 2230
rect 9982 1618 9992 2230
rect 9914 1482 9992 1618
rect 10430 2230 10508 2235
rect 10430 1618 10440 2230
rect 10498 1618 10508 2230
rect 10430 1482 10508 1618
rect 10946 2230 11024 2235
rect 10946 1618 10956 2230
rect 11014 1618 11024 2230
rect 10946 1482 11024 1618
rect 11462 2230 11540 2235
rect 11462 1618 11472 2230
rect 11530 1618 11540 2230
rect 11462 1482 11540 1618
rect 11978 2230 12056 2235
rect 11978 1618 11988 2230
rect 12046 1618 12056 2230
rect 11978 1482 12056 1618
rect 12494 2230 12572 2235
rect 12494 1618 12504 2230
rect 12562 1618 12572 2230
rect 12494 1482 12572 1618
rect 13010 2230 13088 2235
rect 13010 1618 13020 2230
rect 13078 1618 13088 2230
rect 13010 1482 13088 1618
rect 6269 1380 13517 1482
rect 13662 1466 13722 2997
rect 22430 2922 22892 2952
rect 22430 2658 22442 2922
rect 22858 2658 22892 2922
rect 13657 1461 13727 1466
rect 13657 1401 13662 1461
rect 13722 1401 13727 1461
rect 13657 1396 13727 1401
rect 6269 1187 6371 1380
rect 6818 1244 6896 1380
rect 6070 1182 6386 1187
rect 6070 1078 6080 1182
rect 6376 1078 6386 1182
rect 6070 1073 6386 1078
rect 6818 632 6828 1244
rect 6886 632 6896 1244
rect 6818 627 6896 632
rect 7334 1244 7412 1380
rect 7334 632 7344 1244
rect 7402 632 7412 1244
rect 7334 627 7412 632
rect 7850 1244 7928 1380
rect 7850 632 7860 1244
rect 7918 632 7928 1244
rect 7850 627 7928 632
rect 8366 1244 8444 1380
rect 8366 632 8376 1244
rect 8434 632 8444 1244
rect 8366 627 8444 632
rect 8882 1244 8960 1380
rect 8882 632 8892 1244
rect 8950 632 8960 1244
rect 8882 627 8960 632
rect 9398 1244 9476 1380
rect 9398 632 9408 1244
rect 9466 632 9476 1244
rect 9398 627 9476 632
rect 9914 1250 9992 1380
rect 9914 1246 9990 1250
rect 9914 630 9924 1246
rect 9980 630 9990 1246
rect 9914 625 9990 630
rect 10430 1244 10508 1380
rect 10430 632 10440 1244
rect 10498 632 10508 1244
rect 10430 627 10508 632
rect 10946 1244 11024 1380
rect 10946 632 10956 1244
rect 11014 632 11024 1244
rect 10946 627 11024 632
rect 11462 1244 11540 1380
rect 11462 632 11472 1244
rect 11530 632 11540 1244
rect 11462 627 11540 632
rect 11978 1244 12056 1380
rect 11978 632 11988 1244
rect 12046 632 12056 1244
rect 11978 627 12056 632
rect 12494 1244 12572 1380
rect 12494 632 12504 1244
rect 12562 632 12572 1244
rect 12494 627 12572 632
rect 13010 1244 13088 1380
rect 13010 632 13020 1244
rect 13078 632 13088 1244
rect 13010 627 13088 632
rect 13415 98 13517 1380
rect 13415 6 13420 98
rect 13512 6 13517 98
rect 13415 1 13517 6
rect -3750 -588 -3626 -583
rect -3750 -668 -3740 -588
rect -3636 -668 -3626 -588
rect -3750 -673 -3626 -668
rect -4337 -960 -4251 -955
rect -4337 -1036 -4332 -960
rect -4256 -1036 -4251 -960
rect -4337 -1041 -4251 -1036
rect -3722 -1127 -3662 -673
rect -3748 -1132 -3634 -1127
rect -3748 -1208 -3738 -1132
rect -3644 -1208 -3634 -1132
rect -3748 -1213 -3634 -1208
rect -3722 -2259 -3658 -1213
rect -3746 -2264 -3630 -2259
rect -3746 -2356 -3736 -2264
rect -3640 -2356 -3630 -2264
rect -3746 -2361 -3630 -2356
rect -3722 -2813 -3658 -2361
rect -3748 -2818 -3632 -2813
rect -3748 -2910 -3738 -2818
rect -3642 -2910 -3632 -2818
rect -3748 -2915 -3632 -2910
rect 22430 -3592 22892 2658
rect 33426 451 33522 6361
rect 33660 3463 33756 9373
rect 33942 4995 34038 10905
rect 34202 8007 34298 12564
rect 34193 8001 34298 8007
rect 34295 7899 34298 8001
rect 34193 7893 34298 7899
rect 33937 4989 34039 4995
rect 33937 4881 34039 4887
rect 33645 3457 33756 3463
rect 33747 3355 33756 3457
rect 33645 3349 33756 3355
rect 33417 445 33522 451
rect 33519 343 33522 445
rect 33417 337 33522 343
rect 30748 -331 30844 -326
rect 30748 -417 30753 -331
rect 30839 -417 30844 -331
rect 30748 -467 30844 -417
rect 30743 -472 30849 -467
rect 30743 -568 30748 -472
rect 30844 -568 30849 -472
rect 30743 -573 30849 -568
rect 23176 -3592 24032 -3370
rect 22430 -4094 24032 -3592
rect 22430 -4146 22892 -4094
rect 23176 -4212 24032 -4094
rect 33426 -4216 33522 337
rect 33660 -477 33756 3349
rect 33660 -563 33665 -477
rect 33751 -563 33756 -477
rect 33660 -2561 33756 -563
rect 33942 2001 34038 4881
rect 33942 1915 33947 2001
rect 34033 1915 34038 2001
rect 34202 1983 34298 7893
rect 33942 -1029 34038 1915
rect 34197 1977 34299 1983
rect 34197 1869 34299 1875
rect 33933 -1035 34038 -1029
rect 34035 -1137 34038 -1035
rect 33933 -1143 34038 -1137
rect 33653 -2567 33756 -2561
rect 33755 -2669 33756 -2567
rect 33653 -2675 33756 -2669
rect 33660 -4218 33756 -2675
rect 33942 -4208 34038 -1143
rect 34202 1745 34298 1869
rect 34202 1659 34207 1745
rect 34293 1659 34298 1745
rect 34202 -4041 34298 1659
rect 34193 -4047 34298 -4041
rect 34295 -4149 34298 -4047
rect 34193 -4155 34298 -4149
rect 34202 -4226 34298 -4155
<< via3 >>
rect 33423 12391 33525 12493
rect 33941 10911 34043 11013
rect 33653 9379 33755 9481
rect 33417 6367 33519 6469
rect 34193 7899 34295 8001
rect 33937 4887 34039 4989
rect 33645 3355 33747 3457
rect 33417 343 33519 445
rect 34197 1875 34299 1977
rect 33933 -1137 34035 -1035
rect 33653 -2669 33755 -2567
rect 34193 -4149 34295 -4047
<< metal4 >>
rect 33422 12493 34456 12494
rect 33422 12391 33423 12493
rect 33525 12391 34456 12493
rect 33422 12390 34456 12391
rect 33940 11013 34460 11014
rect 33940 10911 33941 11013
rect 34043 10911 34460 11013
rect 33940 10910 34460 10911
rect 33652 9481 34456 9482
rect 33652 9379 33653 9481
rect 33755 9379 34456 9481
rect 33652 9378 34456 9379
rect 34192 8001 34458 8002
rect 34192 7899 34193 8001
rect 34295 7899 34458 8001
rect 34192 7898 34458 7899
rect 33406 6469 34476 6470
rect 33406 6367 33417 6469
rect 33519 6367 34476 6469
rect 33406 6366 34476 6367
rect 33936 4989 34458 4990
rect 33936 4887 33937 4989
rect 34039 4887 34458 4989
rect 33936 4886 34458 4887
rect 33644 3457 34458 3458
rect 33644 3355 33645 3457
rect 33747 3355 34458 3457
rect 33644 3354 34458 3355
rect 34196 1977 34472 1978
rect 34196 1875 34197 1977
rect 34299 1875 34472 1977
rect 34196 1874 34472 1875
rect 33416 445 34456 446
rect 33416 343 33417 445
rect 33519 343 34456 445
rect 33416 342 34456 343
rect 33932 -1035 34484 -1034
rect 33932 -1137 33933 -1035
rect 34035 -1137 34484 -1035
rect 33932 -1138 34484 -1137
rect 33652 -2567 34456 -2566
rect 33652 -2669 33653 -2567
rect 33755 -2669 34456 -2567
rect 33652 -2670 34456 -2669
rect 34192 -4047 34456 -4046
rect 34192 -4149 34193 -4047
rect 34295 -4149 34456 -4047
rect 34192 -4150 34456 -4149
use sky130_fd_pr__cap_mim_m3_1_Z5XS7R  sky130_fd_pr__cap_mim_m3_1_Z5XS7R_1
timestamp 1713452221
transform 0 1 42512 -1 0 4766
box -8916 -8160 8916 8160
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1713465581
transform 1 0 -8469 0 1 3877
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_1
timestamp 1713465581
transform 1 0 -9289 0 1 3883
box -211 -310 211 310
use sky130_fd_pr__nfet_g5v0d10v5_2B7385  sky130_fd_pr__nfet_g5v0d10v5_2B7385_0
timestamp 1713300479
transform 1 0 -579 0 1 558
box -2521 -1058 2521 1058
use sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR  sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR_0
timestamp 1713285936
transform 1 0 27459 0 1 -1342
box -5359 -458 5359 458
use sky130_fd_pr__nfet_g5v0d10v5_79TVLH  sky130_fd_pr__nfet_g5v0d10v5_79TVLH_0
timestamp 1713306471
transform 1 0 9953 0 1 938
box -3553 -558 3553 558
use sky130_fd_pr__nfet_g5v0d10v5_79TVLH  sky130_fd_pr__nfet_g5v0d10v5_79TVLH_1
timestamp 1713306471
transform 1 0 9953 0 1 1924
box -3553 -558 3553 558
use sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z  sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z_0
timestamp 1713297702
transform 1 0 9469 0 1 -592
box -4069 -708 4069 708
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_0
timestamp 1713414983
transform 1 0 -3688 0 1 -900
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_1
timestamp 1713414983
transform 1 0 -3690 0 1 -2588
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_2
timestamp 1713414983
transform 1 0 -1824 0 1 2180
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_3
timestamp 1713414983
transform 1 0 -4764 0 1 -114
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_4
timestamp 1713414983
transform 1 0 -4764 0 1 672
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_5
timestamp 1713414983
transform 1 0 -4764 0 1 1458
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_6
timestamp 1713414983
transform 1 0 -4764 0 1 -900
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_7
timestamp 1713414983
transform 1 0 -4764 0 1 -1686
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_8
timestamp 1713414983
transform 1 0 -4764 0 1 -2472
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_9
timestamp 1713414983
transform 1 0 -4764 0 1 -3258
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_10
timestamp 1713414983
transform 1 0 -5968 0 1 -3262
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_11
timestamp 1713414983
transform 1 0 -5968 0 1 -2476
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_12
timestamp 1713414983
transform 1 0 -5968 0 1 -1690
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_13
timestamp 1713414983
transform 1 0 -5968 0 1 -904
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14
timestamp 1713414983
transform 1 0 -5968 0 1 2240
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_15
timestamp 1713414983
transform 1 0 -5968 0 1 1454
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_16
timestamp 1713414983
transform 1 0 -5968 0 1 668
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_17
timestamp 1713414983
transform 1 0 -5968 0 1 -118
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18
timestamp 1713414983
transform 1 0 -4764 0 1 2244
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_CTEUHA  sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_19
timestamp 1713414983
transform 1 0 -3466 0 1 2180
box -278 -458 278 458
use sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN  sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN_0
timestamp 1713285936
transform 1 0 27211 0 1 -2572
box -5101 -458 5101 458
use sky130_fd_pr__nfet_g5v0d10v5_HG2LSW  sky130_fd_pr__nfet_g5v0d10v5_HG2LSW_0
timestamp 1713291415
transform 1 0 4429 0 1 -2691
box -328 -408 328 408
use sky130_fd_pr__nfet_g5v0d10v5_N64HU4  sky130_fd_pr__nfet_g5v0d10v5_N64HU4_0
timestamp 1713278525
transform 1 0 763 0 1 -1442
box -3863 -458 3863 458
use sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U  sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U_0
timestamp 1713246000
transform 1 0 305 0 1 -2642
box -3405 -458 3405 458
use sky130_fd_pr__nfet_g5v0d10v5_PGZBW9  sky130_fd_pr__nfet_g5v0d10v5_PGZBW9_0
timestamp 1713300419
transform 1 0 17553 0 1 -2242
box -3553 -858 3553 858
use sky130_fd_pr__nfet_g5v0d10v5_RMXH5H  sky130_fd_pr__nfet_g5v0d10v5_RMXH5H_0
timestamp 1713300419
transform 1 0 19847 0 1 1858
box -1747 -458 1747 458
use sky130_fd_pr__nfet_g5v0d10v5_U73S5M  sky130_fd_pr__nfet_g5v0d10v5_U73S5M_0
timestamp 1713300479
transform 1 0 27057 0 1 808
box -4585 -1258 4585 1258
use sky130_fd_pr__nfet_g5v0d10v5_UGZTXE  sky130_fd_pr__nfet_g5v0d10v5_UGZTXE_0
timestamp 1713300419
transform 1 0 17811 0 1 -142
box -3811 -858 3811 858
use sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J  sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J_0
timestamp 1713291448
transform 1 0 9953 0 1 -2392
box -3553 -708 3553 708
use sky130_fd_pr__nfet_g5v0d10v5_USXRNR  sky130_fd_pr__nfet_g5v0d10v5_USXRNR_0
timestamp 1713300419
transform 1 0 15877 0 1 1859
box -1876 -458 1876 458
use sky130_fd_pr__nfet_g5v0d10v5_WK95DB  sky130_fd_pr__nfet_g5v0d10v5_WK95DB_0
timestamp 1713300479
transform 1 0 3489 0 1 208
box -989 -708 989 708
use sky130_fd_pr__nfet_g5v0d10v5_YJ3VXJ  sky130_fd_pr__nfet_g5v0d10v5_YJ3VXJ_0
timestamp 1713416422
transform 1 0 -2645 0 1 2180
box -673 -458 673 458
use sky130_fd_pr__pfet_01v8_U4BBJH  sky130_fd_pr__pfet_01v8_U4BBJH_0
timestamp 1713465581
transform 1 0 -8469 0 1 4612
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_U4BBJH  sky130_fd_pr__pfet_01v8_U4BBJH_1
timestamp 1713465581
transform 1 0 -9289 0 1 4612
box -211 -419 211 419
use sky130_fd_pr__pfet_g5v0d10v5_3QL9S5  sky130_fd_pr__pfet_g5v0d10v5_3QL9S5_0
timestamp 1713408563
transform 1 0 12210 0 1 12285
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_3QL9S5  sky130_fd_pr__pfet_g5v0d10v5_3QL9S5_1
timestamp 1713408563
transform 1 0 13030 0 1 12291
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_AUMBFF  sky130_fd_pr__pfet_g5v0d10v5_AUMBFF_0
timestamp 1713391144
transform 1 0 28313 0 1 6187
box -4615 -2797 4615 2797
use sky130_fd_pr__pfet_g5v0d10v5_BH2H9S  sky130_fd_pr__pfet_g5v0d10v5_BH2H9S_0
timestamp 1713400206
transform 1 0 -327 0 1 10929
box -2551 -1897 2551 1897
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_0
timestamp 1713418706
transform 1 0 1084 0 1 4029
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_1
timestamp 1713418706
transform 1 0 -1204 0 1 7645
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_2
timestamp 1713418706
transform 1 0 1084 0 1 5233
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_3
timestamp 1713418706
transform 1 0 -1204 0 1 6441
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_4
timestamp 1713418706
transform 1 0 -1204 0 1 5237
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_5
timestamp 1713418706
transform 1 0 -3364 0 1 3933
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_6
timestamp 1713418706
transform 1 0 1084 0 1 6437
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_7
timestamp 1713418706
transform 1 0 1084 0 1 7641
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_8
timestamp 1713418706
transform 1 0 124 0 1 5237
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_9
timestamp 1713418706
transform 1 0 124 0 1 4033
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_10
timestamp 1713418706
transform 1 0 124 0 1 7645
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_11
timestamp 1713418706
transform 1 0 124 0 1 6441
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_12
timestamp 1713418706
transform 1 0 -302 0 1 5237
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13
timestamp 1713418706
transform 1 0 -302 0 1 4033
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_14
timestamp 1713418706
transform 1 0 -302 0 1 7645
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_15
timestamp 1713418706
transform 1 0 -302 0 1 6441
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_16
timestamp 1713418706
transform 1 0 -1204 0 1 4033
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_CVG6CD  sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_17
timestamp 1713418706
transform 1 0 -1912 0 1 3945
box -308 -697 308 697
use sky130_fd_pr__pfet_g5v0d10v5_EVM3FM  sky130_fd_pr__pfet_g5v0d10v5_EVM3FM_0
timestamp 1713394428
transform 1 0 10329 0 1 11511
box -1019 -1197 1019 1197
use sky130_fd_pr__pfet_g5v0d10v5_HQ4STX  sky130_fd_pr__pfet_g5v0d10v5_HQ4STX_0
timestamp 1713332554
transform 1 0 23032 0 1 12243
box -358 -597 358 597
use sky130_fd_pr__pfet_g5v0d10v5_PP2RNK  sky130_fd_pr__pfet_g5v0d10v5_PP2RNK_0
timestamp 1713394428
transform 1 0 6155 0 1 8551
box -3325 -1197 3325 1197
use sky130_fd_pr__pfet_g5v0d10v5_Q46EE6  sky130_fd_pr__pfet_g5v0d10v5_Q46EE6_0
timestamp 1713331574
transform 1 0 19671 0 1 12343
box -2035 -497 2035 497
use sky130_fd_pr__pfet_g5v0d10v5_QL2RRT  sky130_fd_pr__pfet_g5v0d10v5_QL2RRT_0
timestamp 1713394428
transform 1 0 6378 0 1 6008
box -3583 -897 3583 897
use sky130_fd_pr__pfet_g5v0d10v5_QL2RRT  sky130_fd_pr__pfet_g5v0d10v5_QL2RRT_1
timestamp 1713394428
transform 1 0 6378 0 1 4404
box -3583 -897 3583 897
use sky130_fd_pr__pfet_g5v0d10v5_QRKB8C  sky130_fd_pr__pfet_g5v0d10v5_QRKB8C_0
timestamp 1713332875
transform 1 0 28455 0 1 12183
box -4873 -697 4873 697
use sky130_fd_pr__pfet_g5v0d10v5_QSKB8C  sky130_fd_pr__pfet_g5v0d10v5_QSKB8C_0
timestamp 1713390278
transform 1 0 27831 0 1 10263
box -5131 -697 5131 697
use sky130_fd_pr__pfet_g5v0d10v5_QTY6H6  sky130_fd_pr__pfet_g5v0d10v5_QTY6H6_0
timestamp 1713331128
transform 1 0 15217 0 1 12357
box -1777 -497 1777 497
use sky130_fd_pr__pfet_g5v0d10v5_QTY6KC  sky130_fd_pr__pfet_g5v0d10v5_QTY6KC_0
timestamp 1713393095
transform 1 0 19983 0 1 4087
box -1777 -697 1777 697
use sky130_fd_pr__pfet_g5v0d10v5_TT9EEV  sky130_fd_pr__pfet_g5v0d10v5_TT9EEV_0
timestamp 1713393126
transform 1 0 15324 0 1 4071
box -1906 -717 1906 717
use sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD  sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD_1
timestamp 1713416651
transform 1 0 -2649 0 1 5343
box -1019 -697 1019 697
use sky130_fd_pr__pfet_g5v0d10v5_W75H7K  sky130_fd_pr__pfet_g5v0d10v5_W75H7K_0
timestamp 1713394428
transform 1 0 16891 0 1 9933
box -5131 -1497 5131 1497
use sky130_fd_pr__pfet_g5v0d10v5_WKXP7K  sky130_fd_pr__pfet_g5v0d10v5_WKXP7K_0
timestamp 1713393625
transform 1 0 16649 0 1 6651
box -5389 -1497 5389 1497
use sky130_fd_pr__pfet_g5v0d10v5_XW23Q2  sky130_fd_pr__pfet_g5v0d10v5_XW23Q2_0
timestamp 1713394428
transform 1 0 5909 0 1 11511
box -3067 -1197 3067 1197
use sky130_fd_pr__res_generic_po_U7N8A7  sky130_fd_pr__res_generic_po_U7N8A7_0
timestamp 1713451382
transform 1 0 32463 0 1 644
box -755 -1096 755 1096
<< labels >>
flabel metal2 -4352 5632 -3966 6052 0 FreeSans 960 0 0 0 vinn
port 4 nsew
flabel metal2 -4352 6252 -3966 6672 0 FreeSans 960 0 0 0 vinp
port 5 nsew
flabel metal2 -4344 6842 -3958 7262 0 FreeSans 960 0 0 0 ibias
port 3 nsew
flabel metal3 23214 -4164 23930 -3444 0 FreeSans 1920 0 0 0 vout
port 2 nsew
flabel metal1 -6048 -5544 -4866 -4798 0 FreeSans 3200 0 0 0 avss
port 6 nsew
flabel metal1 -5166 14382 -3852 15374 0 FreeSans 3200 0 0 0 avdd
port 1 nsew
flabel viali -9940 3461 -9572 3611 0 FreeSans 640 0 0 0 dvss
port 8 nsew
flabel viali -9948 4991 -9580 5141 0 FreeSans 640 0 0 0 dvdd
port 7 nsew
flabel metal1 -9950 4095 -9694 4363 0 FreeSans 640 0 0 0 ena
port 9 nsew
flabel locali 6836 -3118 6962 -3090 0 FreeSans 640 0 0 0 vb4
flabel metal2 5524 -1118 5598 -1070 0 FreeSans 480 0 0 0 vb3
flabel metal1 6232 -1256 6334 -1224 0 FreeSans 320 0 0 0 net28
flabel metal1 7802 -1248 7904 -1216 0 FreeSans 320 0 0 0 net29
flabel metal1 11712 -1248 11810 -1226 0 FreeSans 320 0 0 0 net12
flabel metal1 27878 -1730 27930 -1712 0 FreeSans 320 0 0 0 net16
flabel metal1 24832 -1720 24832 -1720 0 FreeSans 320 0 0 0 net24
flabel metal2 21926 -886 22036 -850 0 FreeSans 320 0 0 0 vb7
flabel metal1 22922 -2482 22922 -2482 0 FreeSans 320 0 0 0 vb8
flabel metal1 31010 -1734 31096 -1714 0 FreeSans 320 0 0 0 net25
flabel metal2 -1124 -3262 -1124 -3262 0 FreeSans 320 0 0 0 net31
flabel metal2 -3100 -3102 -3100 -3102 0 FreeSans 320 0 0 0 net34
flabel metal2 -150 -2226 -150 -2226 0 FreeSans 320 0 0 0 net20
flabel metal2 18178 11510 18178 11510 0 FreeSans 320 0 0 0 net21
flabel metal2 18028 12744 18028 12744 0 FreeSans 320 0 0 0 net32
flabel metal1 14774 11950 14774 11950 0 FreeSans 320 0 0 0 net22
flabel metal2 -1588 -856 -1034 -826 0 FreeSans 320 0 0 0 net33
flabel metal3 6288 1396 6288 1396 0 FreeSans 320 0 0 0 vtailn
flabel metal3 9760 5184 9760 5184 0 FreeSans 320 0 0 0 vtailp
flabel metal2 27138 11700 27138 11700 0 FreeSans 320 0 0 0 vb5
flabel metal2 27024 9786 27024 9786 0 FreeSans 320 0 0 0 vb6
flabel metal2 15820 11176 15820 11176 0 FreeSans 320 0 0 0 net5
flabel metal2 15060 7886 15060 7886 0 FreeSans 320 0 0 0 vb2
flabel metal1 13656 8032 13656 8032 0 FreeSans 320 0 0 0 net3
flabel metal1 18714 8030 18714 8030 0 FreeSans 320 0 0 0 net4
flabel metal2 17550 -812 17550 -812 0 FreeSans 320 0 0 0 vb3
flabel metal1 -2820 1812 -2820 1812 0 FreeSans 320 0 0 0 net35
flabel metal1 3470 850 3470 850 0 FreeSans 320 0 0 0 net18
flabel metal1 7914 24 7914 24 0 FreeSans 320 0 0 0 vb1
flabel metal1 15154 1442 15154 1442 0 FreeSans 320 0 0 0 net6
flabel metal1 18928 2190 18928 2190 0 FreeSans 320 0 0 0 net10
flabel metal1 16744 1452 16744 1452 0 FreeSans 320 0 0 0 net8
flabel metal1 29586 9676 29586 9676 0 FreeSans 320 0 0 0 net10
flabel metal1 29606 10844 29606 10844 0 FreeSans 320 0 0 0 net13
flabel metal1 -3628 3170 -3628 3170 0 FreeSans 320 0 0 0 enab_avdd
flabel metal2 17372 -1422 17372 -1422 0 FreeSans 320 0 0 0 net1
flabel metal1 19564 -1108 19564 -1108 0 FreeSans 320 0 0 0 net2
flabel metal2 -2646 12570 -2646 12576 0 FreeSans 320 0 0 0 net18
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713394428
<< error_p >>
rect -743 981 -679 987
rect -585 981 -521 987
rect -427 981 -363 987
rect -269 981 -205 987
rect -111 981 -47 987
rect 47 981 111 987
rect 205 981 269 987
rect 363 981 427 987
rect 521 981 585 987
rect 679 981 743 987
rect -743 947 -731 981
rect -585 947 -573 981
rect -427 947 -415 981
rect -269 947 -257 981
rect -111 947 -99 981
rect 47 947 59 981
rect 205 947 217 981
rect 363 947 375 981
rect 521 947 533 981
rect 679 947 691 981
rect -743 941 -679 947
rect -585 941 -521 947
rect -427 941 -363 947
rect -269 941 -205 947
rect -111 941 -47 947
rect 47 941 111 947
rect 205 941 269 947
rect 363 941 427 947
rect 521 941 585 947
rect 679 941 743 947
rect -743 -947 -679 -941
rect -585 -947 -521 -941
rect -427 -947 -363 -941
rect -269 -947 -205 -941
rect -111 -947 -47 -941
rect 47 -947 111 -941
rect 205 -947 269 -941
rect 363 -947 427 -941
rect 521 -947 585 -941
rect 679 -947 743 -941
rect -743 -981 -731 -947
rect -585 -981 -573 -947
rect -427 -981 -415 -947
rect -269 -981 -257 -947
rect -111 -981 -99 -947
rect 47 -981 59 -947
rect 205 -981 217 -947
rect 363 -981 375 -947
rect 521 -981 533 -947
rect 679 -981 691 -947
rect -743 -987 -679 -981
rect -585 -987 -521 -981
rect -427 -987 -363 -981
rect -269 -987 -205 -981
rect -111 -987 -47 -981
rect 47 -987 111 -981
rect 205 -987 269 -981
rect 363 -987 427 -981
rect 521 -987 585 -981
rect 679 -987 743 -981
<< nwell >>
rect -1019 -1197 1019 1197
<< mvpmos >>
rect -761 -900 -661 900
rect -603 -900 -503 900
rect -445 -900 -345 900
rect -287 -900 -187 900
rect -129 -900 -29 900
rect 29 -900 129 900
rect 187 -900 287 900
rect 345 -900 445 900
rect 503 -900 603 900
rect 661 -900 761 900
<< mvpdiff >>
rect -819 888 -761 900
rect -819 -888 -807 888
rect -773 -888 -761 888
rect -819 -900 -761 -888
rect -661 888 -603 900
rect -661 -888 -649 888
rect -615 -888 -603 888
rect -661 -900 -603 -888
rect -503 888 -445 900
rect -503 -888 -491 888
rect -457 -888 -445 888
rect -503 -900 -445 -888
rect -345 888 -287 900
rect -345 -888 -333 888
rect -299 -888 -287 888
rect -345 -900 -287 -888
rect -187 888 -129 900
rect -187 -888 -175 888
rect -141 -888 -129 888
rect -187 -900 -129 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 129 888 187 900
rect 129 -888 141 888
rect 175 -888 187 888
rect 129 -900 187 -888
rect 287 888 345 900
rect 287 -888 299 888
rect 333 -888 345 888
rect 287 -900 345 -888
rect 445 888 503 900
rect 445 -888 457 888
rect 491 -888 503 888
rect 445 -900 503 -888
rect 603 888 661 900
rect 603 -888 615 888
rect 649 -888 661 888
rect 603 -900 661 -888
rect 761 888 819 900
rect 761 -888 773 888
rect 807 -888 819 888
rect 761 -900 819 -888
<< mvpdiffc >>
rect -807 -888 -773 888
rect -649 -888 -615 888
rect -491 -888 -457 888
rect -333 -888 -299 888
rect -175 -888 -141 888
rect -17 -888 17 888
rect 141 -888 175 888
rect 299 -888 333 888
rect 457 -888 491 888
rect 615 -888 649 888
rect 773 -888 807 888
<< mvnsubdiff >>
rect -953 1119 953 1131
rect -953 1085 -845 1119
rect 845 1085 953 1119
rect -953 1073 953 1085
rect -953 1023 -895 1073
rect -953 -1023 -941 1023
rect -907 -1023 -895 1023
rect 895 1023 953 1073
rect -953 -1073 -895 -1023
rect 895 -1023 907 1023
rect 941 -1023 953 1023
rect 895 -1073 953 -1023
rect -953 -1085 953 -1073
rect -953 -1119 -845 -1085
rect 845 -1119 953 -1085
rect -953 -1131 953 -1119
<< mvnsubdiffcont >>
rect -845 1085 845 1119
rect -941 -1023 -907 1023
rect 907 -1023 941 1023
rect -845 -1119 845 -1085
<< poly >>
rect -747 981 -675 997
rect -747 964 -731 981
rect -761 947 -731 964
rect -691 964 -675 981
rect -589 981 -517 997
rect -589 964 -573 981
rect -691 947 -661 964
rect -761 900 -661 947
rect -603 947 -573 964
rect -533 964 -517 981
rect -431 981 -359 997
rect -431 964 -415 981
rect -533 947 -503 964
rect -603 900 -503 947
rect -445 947 -415 964
rect -375 964 -359 981
rect -273 981 -201 997
rect -273 964 -257 981
rect -375 947 -345 964
rect -445 900 -345 947
rect -287 947 -257 964
rect -217 964 -201 981
rect -115 981 -43 997
rect -115 964 -99 981
rect -217 947 -187 964
rect -287 900 -187 947
rect -129 947 -99 964
rect -59 964 -43 981
rect 43 981 115 997
rect 43 964 59 981
rect -59 947 -29 964
rect -129 900 -29 947
rect 29 947 59 964
rect 99 964 115 981
rect 201 981 273 997
rect 201 964 217 981
rect 99 947 129 964
rect 29 900 129 947
rect 187 947 217 964
rect 257 964 273 981
rect 359 981 431 997
rect 359 964 375 981
rect 257 947 287 964
rect 187 900 287 947
rect 345 947 375 964
rect 415 964 431 981
rect 517 981 589 997
rect 517 964 533 981
rect 415 947 445 964
rect 345 900 445 947
rect 503 947 533 964
rect 573 964 589 981
rect 675 981 747 997
rect 675 964 691 981
rect 573 947 603 964
rect 503 900 603 947
rect 661 947 691 964
rect 731 964 747 981
rect 731 947 761 964
rect 661 900 761 947
rect -761 -947 -661 -900
rect -761 -964 -731 -947
rect -747 -981 -731 -964
rect -691 -964 -661 -947
rect -603 -947 -503 -900
rect -603 -964 -573 -947
rect -691 -981 -675 -964
rect -747 -997 -675 -981
rect -589 -981 -573 -964
rect -533 -964 -503 -947
rect -445 -947 -345 -900
rect -445 -964 -415 -947
rect -533 -981 -517 -964
rect -589 -997 -517 -981
rect -431 -981 -415 -964
rect -375 -964 -345 -947
rect -287 -947 -187 -900
rect -287 -964 -257 -947
rect -375 -981 -359 -964
rect -431 -997 -359 -981
rect -273 -981 -257 -964
rect -217 -964 -187 -947
rect -129 -947 -29 -900
rect -129 -964 -99 -947
rect -217 -981 -201 -964
rect -273 -997 -201 -981
rect -115 -981 -99 -964
rect -59 -964 -29 -947
rect 29 -947 129 -900
rect 29 -964 59 -947
rect -59 -981 -43 -964
rect -115 -997 -43 -981
rect 43 -981 59 -964
rect 99 -964 129 -947
rect 187 -947 287 -900
rect 187 -964 217 -947
rect 99 -981 115 -964
rect 43 -997 115 -981
rect 201 -981 217 -964
rect 257 -964 287 -947
rect 345 -947 445 -900
rect 345 -964 375 -947
rect 257 -981 273 -964
rect 201 -997 273 -981
rect 359 -981 375 -964
rect 415 -964 445 -947
rect 503 -947 603 -900
rect 503 -964 533 -947
rect 415 -981 431 -964
rect 359 -997 431 -981
rect 517 -981 533 -964
rect 573 -964 603 -947
rect 661 -947 761 -900
rect 661 -964 691 -947
rect 573 -981 589 -964
rect 517 -997 589 -981
rect 675 -981 691 -964
rect 731 -964 761 -947
rect 731 -981 747 -964
rect 675 -997 747 -981
<< polycont >>
rect -731 947 -691 981
rect -573 947 -533 981
rect -415 947 -375 981
rect -257 947 -217 981
rect -99 947 -59 981
rect 59 947 99 981
rect 217 947 257 981
rect 375 947 415 981
rect 533 947 573 981
rect 691 947 731 981
rect -731 -981 -691 -947
rect -573 -981 -533 -947
rect -415 -981 -375 -947
rect -257 -981 -217 -947
rect -99 -981 -59 -947
rect 59 -981 99 -947
rect 217 -981 257 -947
rect 375 -981 415 -947
rect 533 -981 573 -947
rect 691 -981 731 -947
<< locali >>
rect -941 1085 -845 1119
rect 845 1085 941 1119
rect -941 1023 -907 1085
rect 907 1023 941 1085
rect -747 947 -731 981
rect -691 947 -675 981
rect -589 947 -573 981
rect -533 947 -517 981
rect -431 947 -415 981
rect -375 947 -359 981
rect -273 947 -257 981
rect -217 947 -201 981
rect -115 947 -99 981
rect -59 947 -43 981
rect 43 947 59 981
rect 99 947 115 981
rect 201 947 217 981
rect 257 947 273 981
rect 359 947 375 981
rect 415 947 431 981
rect 517 947 533 981
rect 573 947 589 981
rect 675 947 691 981
rect 731 947 747 981
rect -807 888 -773 904
rect -807 -904 -773 -888
rect -649 888 -615 904
rect -649 -904 -615 -888
rect -491 888 -457 904
rect -491 -904 -457 -888
rect -333 888 -299 904
rect -333 -904 -299 -888
rect -175 888 -141 904
rect -175 -904 -141 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 141 888 175 904
rect 141 -904 175 -888
rect 299 888 333 904
rect 299 -904 333 -888
rect 457 888 491 904
rect 457 -904 491 -888
rect 615 888 649 904
rect 615 -904 649 -888
rect 773 888 807 904
rect 773 -904 807 -888
rect -747 -981 -731 -947
rect -691 -981 -675 -947
rect -589 -981 -573 -947
rect -533 -981 -517 -947
rect -431 -981 -415 -947
rect -375 -981 -359 -947
rect -273 -981 -257 -947
rect -217 -981 -201 -947
rect -115 -981 -99 -947
rect -59 -981 -43 -947
rect 43 -981 59 -947
rect 99 -981 115 -947
rect 201 -981 217 -947
rect 257 -981 273 -947
rect 359 -981 375 -947
rect 415 -981 431 -947
rect 517 -981 533 -947
rect 573 -981 589 -947
rect 675 -981 691 -947
rect 731 -981 747 -947
rect -941 -1085 -907 -1023
rect 907 -1085 941 -1023
rect -941 -1119 -845 -1085
rect 845 -1119 941 -1085
<< viali >>
rect -731 947 -691 981
rect -573 947 -533 981
rect -415 947 -375 981
rect -257 947 -217 981
rect -99 947 -59 981
rect 59 947 99 981
rect 217 947 257 981
rect 375 947 415 981
rect 533 947 573 981
rect 691 947 731 981
rect -807 -888 -773 888
rect -649 -888 -615 888
rect -491 -888 -457 888
rect -333 -888 -299 888
rect -175 -888 -141 888
rect -17 -888 17 888
rect 141 -888 175 888
rect 299 -888 333 888
rect 457 -888 491 888
rect 615 -888 649 888
rect 773 -888 807 888
rect -731 -981 -691 -947
rect -573 -981 -533 -947
rect -415 -981 -375 -947
rect -257 -981 -217 -947
rect -99 -981 -59 -947
rect 59 -981 99 -947
rect 217 -981 257 -947
rect 375 -981 415 -947
rect 533 -981 573 -947
rect 691 -981 731 -947
<< metal1 >>
rect -743 981 -679 987
rect -743 947 -731 981
rect -691 947 -679 981
rect -743 941 -679 947
rect -585 981 -521 987
rect -585 947 -573 981
rect -533 947 -521 981
rect -585 941 -521 947
rect -427 981 -363 987
rect -427 947 -415 981
rect -375 947 -363 981
rect -427 941 -363 947
rect -269 981 -205 987
rect -269 947 -257 981
rect -217 947 -205 981
rect -269 941 -205 947
rect -111 981 -47 987
rect -111 947 -99 981
rect -59 947 -47 981
rect -111 941 -47 947
rect 47 981 111 987
rect 47 947 59 981
rect 99 947 111 981
rect 47 941 111 947
rect 205 981 269 987
rect 205 947 217 981
rect 257 947 269 981
rect 205 941 269 947
rect 363 981 427 987
rect 363 947 375 981
rect 415 947 427 981
rect 363 941 427 947
rect 521 981 585 987
rect 521 947 533 981
rect 573 947 585 981
rect 521 941 585 947
rect 679 981 743 987
rect 679 947 691 981
rect 731 947 743 981
rect 679 941 743 947
rect -813 888 -767 900
rect -813 -888 -807 888
rect -773 -888 -767 888
rect -813 -900 -767 -888
rect -655 888 -609 900
rect -655 -888 -649 888
rect -615 -888 -609 888
rect -655 -900 -609 -888
rect -497 888 -451 900
rect -497 -888 -491 888
rect -457 -888 -451 888
rect -497 -900 -451 -888
rect -339 888 -293 900
rect -339 -888 -333 888
rect -299 -888 -293 888
rect -339 -900 -293 -888
rect -181 888 -135 900
rect -181 -888 -175 888
rect -141 -888 -135 888
rect -181 -900 -135 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 135 888 181 900
rect 135 -888 141 888
rect 175 -888 181 888
rect 135 -900 181 -888
rect 293 888 339 900
rect 293 -888 299 888
rect 333 -888 339 888
rect 293 -900 339 -888
rect 451 888 497 900
rect 451 -888 457 888
rect 491 -888 497 888
rect 451 -900 497 -888
rect 609 888 655 900
rect 609 -888 615 888
rect 649 -888 655 888
rect 609 -900 655 -888
rect 767 888 813 900
rect 767 -888 773 888
rect 807 -888 813 888
rect 767 -900 813 -888
rect -743 -947 -679 -941
rect -743 -981 -731 -947
rect -691 -981 -679 -947
rect -743 -987 -679 -981
rect -585 -947 -521 -941
rect -585 -981 -573 -947
rect -533 -981 -521 -947
rect -585 -987 -521 -981
rect -427 -947 -363 -941
rect -427 -981 -415 -947
rect -375 -981 -363 -947
rect -427 -987 -363 -981
rect -269 -947 -205 -941
rect -269 -981 -257 -947
rect -217 -981 -205 -947
rect -269 -987 -205 -981
rect -111 -947 -47 -941
rect -111 -981 -99 -947
rect -59 -981 -47 -947
rect -111 -987 -47 -981
rect 47 -947 111 -941
rect 47 -981 59 -947
rect 99 -981 111 -947
rect 47 -987 111 -981
rect 205 -947 269 -941
rect 205 -981 217 -947
rect 257 -981 269 -947
rect 205 -987 269 -981
rect 363 -947 427 -941
rect 363 -981 375 -947
rect 415 -981 427 -947
rect 363 -987 427 -981
rect 521 -947 585 -941
rect 521 -981 533 -947
rect 573 -981 585 -947
rect 521 -987 585 -981
rect 679 -947 743 -941
rect 679 -981 691 -947
rect 731 -981 743 -947
rect 679 -987 743 -981
<< properties >>
string FIXED_BBOX -924 -1102 924 1102
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9 l 0.5 m 1 nf 10 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

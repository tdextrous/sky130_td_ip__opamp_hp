magic
tech sky130A
magscale 1 2
timestamp 1713278525
<< pwell >>
rect -3863 -458 3863 458
<< mvnmos >>
rect -3635 -200 -3235 200
rect -3177 -200 -2777 200
rect -2719 -200 -2319 200
rect -2261 -200 -1861 200
rect -1803 -200 -1403 200
rect -1345 -200 -945 200
rect -887 -200 -487 200
rect -429 -200 -29 200
rect 29 -200 429 200
rect 487 -200 887 200
rect 945 -200 1345 200
rect 1403 -200 1803 200
rect 1861 -200 2261 200
rect 2319 -200 2719 200
rect 2777 -200 3177 200
rect 3235 -200 3635 200
<< mvndiff >>
rect -3693 188 -3635 200
rect -3693 -188 -3681 188
rect -3647 -188 -3635 188
rect -3693 -200 -3635 -188
rect -3235 188 -3177 200
rect -3235 -188 -3223 188
rect -3189 -188 -3177 188
rect -3235 -200 -3177 -188
rect -2777 188 -2719 200
rect -2777 -188 -2765 188
rect -2731 -188 -2719 188
rect -2777 -200 -2719 -188
rect -2319 188 -2261 200
rect -2319 -188 -2307 188
rect -2273 -188 -2261 188
rect -2319 -200 -2261 -188
rect -1861 188 -1803 200
rect -1861 -188 -1849 188
rect -1815 -188 -1803 188
rect -1861 -200 -1803 -188
rect -1403 188 -1345 200
rect -1403 -188 -1391 188
rect -1357 -188 -1345 188
rect -1403 -200 -1345 -188
rect -945 188 -887 200
rect -945 -188 -933 188
rect -899 -188 -887 188
rect -945 -200 -887 -188
rect -487 188 -429 200
rect -487 -188 -475 188
rect -441 -188 -429 188
rect -487 -200 -429 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 429 188 487 200
rect 429 -188 441 188
rect 475 -188 487 188
rect 429 -200 487 -188
rect 887 188 945 200
rect 887 -188 899 188
rect 933 -188 945 188
rect 887 -200 945 -188
rect 1345 188 1403 200
rect 1345 -188 1357 188
rect 1391 -188 1403 188
rect 1345 -200 1403 -188
rect 1803 188 1861 200
rect 1803 -188 1815 188
rect 1849 -188 1861 188
rect 1803 -200 1861 -188
rect 2261 188 2319 200
rect 2261 -188 2273 188
rect 2307 -188 2319 188
rect 2261 -200 2319 -188
rect 2719 188 2777 200
rect 2719 -188 2731 188
rect 2765 -188 2777 188
rect 2719 -200 2777 -188
rect 3177 188 3235 200
rect 3177 -188 3189 188
rect 3223 -188 3235 188
rect 3177 -200 3235 -188
rect 3635 188 3693 200
rect 3635 -188 3647 188
rect 3681 -188 3693 188
rect 3635 -200 3693 -188
<< mvndiffc >>
rect -3681 -188 -3647 188
rect -3223 -188 -3189 188
rect -2765 -188 -2731 188
rect -2307 -188 -2273 188
rect -1849 -188 -1815 188
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect 1815 -188 1849 188
rect 2273 -188 2307 188
rect 2731 -188 2765 188
rect 3189 -188 3223 188
rect 3647 -188 3681 188
<< mvpsubdiff >>
rect -3827 410 3827 422
rect -3827 376 -3719 410
rect 3719 376 3827 410
rect -3827 364 3827 376
rect -3827 314 -3769 364
rect -3827 -314 -3815 314
rect -3781 -314 -3769 314
rect 3769 314 3827 364
rect -3827 -364 -3769 -314
rect 3769 -314 3781 314
rect 3815 -314 3827 314
rect 3769 -364 3827 -314
rect -3827 -376 3827 -364
rect -3827 -410 -3719 -376
rect 3719 -410 3827 -376
rect -3827 -422 3827 -410
<< mvpsubdiffcont >>
rect -3719 376 3719 410
rect -3815 -314 -3781 314
rect 3781 -314 3815 314
rect -3719 -410 3719 -376
<< poly >>
rect -3561 272 -3309 288
rect -3561 255 -3545 272
rect -3635 238 -3545 255
rect -3325 255 -3309 272
rect -3103 272 -2851 288
rect -3103 255 -3087 272
rect -3325 238 -3235 255
rect -3635 200 -3235 238
rect -3177 238 -3087 255
rect -2867 255 -2851 272
rect -2645 272 -2393 288
rect -2645 255 -2629 272
rect -2867 238 -2777 255
rect -3177 200 -2777 238
rect -2719 238 -2629 255
rect -2409 255 -2393 272
rect -2187 272 -1935 288
rect -2187 255 -2171 272
rect -2409 238 -2319 255
rect -2719 200 -2319 238
rect -2261 238 -2171 255
rect -1951 255 -1935 272
rect -1729 272 -1477 288
rect -1729 255 -1713 272
rect -1951 238 -1861 255
rect -2261 200 -1861 238
rect -1803 238 -1713 255
rect -1493 255 -1477 272
rect -1271 272 -1019 288
rect -1271 255 -1255 272
rect -1493 238 -1403 255
rect -1803 200 -1403 238
rect -1345 238 -1255 255
rect -1035 255 -1019 272
rect -813 272 -561 288
rect -813 255 -797 272
rect -1035 238 -945 255
rect -1345 200 -945 238
rect -887 238 -797 255
rect -577 255 -561 272
rect -355 272 -103 288
rect -355 255 -339 272
rect -577 238 -487 255
rect -887 200 -487 238
rect -429 238 -339 255
rect -119 255 -103 272
rect 103 272 355 288
rect 103 255 119 272
rect -119 238 -29 255
rect -429 200 -29 238
rect 29 238 119 255
rect 339 255 355 272
rect 561 272 813 288
rect 561 255 577 272
rect 339 238 429 255
rect 29 200 429 238
rect 487 238 577 255
rect 797 255 813 272
rect 1019 272 1271 288
rect 1019 255 1035 272
rect 797 238 887 255
rect 487 200 887 238
rect 945 238 1035 255
rect 1255 255 1271 272
rect 1477 272 1729 288
rect 1477 255 1493 272
rect 1255 238 1345 255
rect 945 200 1345 238
rect 1403 238 1493 255
rect 1713 255 1729 272
rect 1935 272 2187 288
rect 1935 255 1951 272
rect 1713 238 1803 255
rect 1403 200 1803 238
rect 1861 238 1951 255
rect 2171 255 2187 272
rect 2393 272 2645 288
rect 2393 255 2409 272
rect 2171 238 2261 255
rect 1861 200 2261 238
rect 2319 238 2409 255
rect 2629 255 2645 272
rect 2851 272 3103 288
rect 2851 255 2867 272
rect 2629 238 2719 255
rect 2319 200 2719 238
rect 2777 238 2867 255
rect 3087 255 3103 272
rect 3309 272 3561 288
rect 3309 255 3325 272
rect 3087 238 3177 255
rect 2777 200 3177 238
rect 3235 238 3325 255
rect 3545 255 3561 272
rect 3545 238 3635 255
rect 3235 200 3635 238
rect -3635 -238 -3235 -200
rect -3635 -255 -3545 -238
rect -3561 -272 -3545 -255
rect -3325 -255 -3235 -238
rect -3177 -238 -2777 -200
rect -3177 -255 -3087 -238
rect -3325 -272 -3309 -255
rect -3561 -288 -3309 -272
rect -3103 -272 -3087 -255
rect -2867 -255 -2777 -238
rect -2719 -238 -2319 -200
rect -2719 -255 -2629 -238
rect -2867 -272 -2851 -255
rect -3103 -288 -2851 -272
rect -2645 -272 -2629 -255
rect -2409 -255 -2319 -238
rect -2261 -238 -1861 -200
rect -2261 -255 -2171 -238
rect -2409 -272 -2393 -255
rect -2645 -288 -2393 -272
rect -2187 -272 -2171 -255
rect -1951 -255 -1861 -238
rect -1803 -238 -1403 -200
rect -1803 -255 -1713 -238
rect -1951 -272 -1935 -255
rect -2187 -288 -1935 -272
rect -1729 -272 -1713 -255
rect -1493 -255 -1403 -238
rect -1345 -238 -945 -200
rect -1345 -255 -1255 -238
rect -1493 -272 -1477 -255
rect -1729 -288 -1477 -272
rect -1271 -272 -1255 -255
rect -1035 -255 -945 -238
rect -887 -238 -487 -200
rect -887 -255 -797 -238
rect -1035 -272 -1019 -255
rect -1271 -288 -1019 -272
rect -813 -272 -797 -255
rect -577 -255 -487 -238
rect -429 -238 -29 -200
rect -429 -255 -339 -238
rect -577 -272 -561 -255
rect -813 -288 -561 -272
rect -355 -272 -339 -255
rect -119 -255 -29 -238
rect 29 -238 429 -200
rect 29 -255 119 -238
rect -119 -272 -103 -255
rect -355 -288 -103 -272
rect 103 -272 119 -255
rect 339 -255 429 -238
rect 487 -238 887 -200
rect 487 -255 577 -238
rect 339 -272 355 -255
rect 103 -288 355 -272
rect 561 -272 577 -255
rect 797 -255 887 -238
rect 945 -238 1345 -200
rect 945 -255 1035 -238
rect 797 -272 813 -255
rect 561 -288 813 -272
rect 1019 -272 1035 -255
rect 1255 -255 1345 -238
rect 1403 -238 1803 -200
rect 1403 -255 1493 -238
rect 1255 -272 1271 -255
rect 1019 -288 1271 -272
rect 1477 -272 1493 -255
rect 1713 -255 1803 -238
rect 1861 -238 2261 -200
rect 1861 -255 1951 -238
rect 1713 -272 1729 -255
rect 1477 -288 1729 -272
rect 1935 -272 1951 -255
rect 2171 -255 2261 -238
rect 2319 -238 2719 -200
rect 2319 -255 2409 -238
rect 2171 -272 2187 -255
rect 1935 -288 2187 -272
rect 2393 -272 2409 -255
rect 2629 -255 2719 -238
rect 2777 -238 3177 -200
rect 2777 -255 2867 -238
rect 2629 -272 2645 -255
rect 2393 -288 2645 -272
rect 2851 -272 2867 -255
rect 3087 -255 3177 -238
rect 3235 -238 3635 -200
rect 3235 -255 3325 -238
rect 3087 -272 3103 -255
rect 2851 -288 3103 -272
rect 3309 -272 3325 -255
rect 3545 -255 3635 -238
rect 3545 -272 3561 -255
rect 3309 -288 3561 -272
<< polycont >>
rect -3545 238 -3325 272
rect -3087 238 -2867 272
rect -2629 238 -2409 272
rect -2171 238 -1951 272
rect -1713 238 -1493 272
rect -1255 238 -1035 272
rect -797 238 -577 272
rect -339 238 -119 272
rect 119 238 339 272
rect 577 238 797 272
rect 1035 238 1255 272
rect 1493 238 1713 272
rect 1951 238 2171 272
rect 2409 238 2629 272
rect 2867 238 3087 272
rect 3325 238 3545 272
rect -3545 -272 -3325 -238
rect -3087 -272 -2867 -238
rect -2629 -272 -2409 -238
rect -2171 -272 -1951 -238
rect -1713 -272 -1493 -238
rect -1255 -272 -1035 -238
rect -797 -272 -577 -238
rect -339 -272 -119 -238
rect 119 -272 339 -238
rect 577 -272 797 -238
rect 1035 -272 1255 -238
rect 1493 -272 1713 -238
rect 1951 -272 2171 -238
rect 2409 -272 2629 -238
rect 2867 -272 3087 -238
rect 3325 -272 3545 -238
<< locali >>
rect -3815 376 -3719 410
rect 3719 376 3815 410
rect -3815 314 -3781 376
rect 3781 314 3815 376
rect -3561 238 -3545 272
rect -3325 238 -3309 272
rect -3103 238 -3087 272
rect -2867 238 -2851 272
rect -2645 238 -2629 272
rect -2409 238 -2393 272
rect -2187 238 -2171 272
rect -1951 238 -1935 272
rect -1729 238 -1713 272
rect -1493 238 -1477 272
rect -1271 238 -1255 272
rect -1035 238 -1019 272
rect -813 238 -797 272
rect -577 238 -561 272
rect -355 238 -339 272
rect -119 238 -103 272
rect 103 238 119 272
rect 339 238 355 272
rect 561 238 577 272
rect 797 238 813 272
rect 1019 238 1035 272
rect 1255 238 1271 272
rect 1477 238 1493 272
rect 1713 238 1729 272
rect 1935 238 1951 272
rect 2171 238 2187 272
rect 2393 238 2409 272
rect 2629 238 2645 272
rect 2851 238 2867 272
rect 3087 238 3103 272
rect 3309 238 3325 272
rect 3545 238 3561 272
rect -3681 188 -3647 204
rect -3681 -204 -3647 -188
rect -3223 188 -3189 204
rect -3223 -204 -3189 -188
rect -2765 188 -2731 204
rect -2765 -204 -2731 -188
rect -2307 188 -2273 204
rect -2307 -204 -2273 -188
rect -1849 188 -1815 204
rect -1849 -204 -1815 -188
rect -1391 188 -1357 204
rect -1391 -204 -1357 -188
rect -933 188 -899 204
rect -933 -204 -899 -188
rect -475 188 -441 204
rect -475 -204 -441 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 441 188 475 204
rect 441 -204 475 -188
rect 899 188 933 204
rect 899 -204 933 -188
rect 1357 188 1391 204
rect 1357 -204 1391 -188
rect 1815 188 1849 204
rect 1815 -204 1849 -188
rect 2273 188 2307 204
rect 2273 -204 2307 -188
rect 2731 188 2765 204
rect 2731 -204 2765 -188
rect 3189 188 3223 204
rect 3189 -204 3223 -188
rect 3647 188 3681 204
rect 3647 -204 3681 -188
rect -3561 -272 -3545 -238
rect -3325 -272 -3309 -238
rect -3103 -272 -3087 -238
rect -2867 -272 -2851 -238
rect -2645 -272 -2629 -238
rect -2409 -272 -2393 -238
rect -2187 -272 -2171 -238
rect -1951 -272 -1935 -238
rect -1729 -272 -1713 -238
rect -1493 -272 -1477 -238
rect -1271 -272 -1255 -238
rect -1035 -272 -1019 -238
rect -813 -272 -797 -238
rect -577 -272 -561 -238
rect -355 -272 -339 -238
rect -119 -272 -103 -238
rect 103 -272 119 -238
rect 339 -272 355 -238
rect 561 -272 577 -238
rect 797 -272 813 -238
rect 1019 -272 1035 -238
rect 1255 -272 1271 -238
rect 1477 -272 1493 -238
rect 1713 -272 1729 -238
rect 1935 -272 1951 -238
rect 2171 -272 2187 -238
rect 2393 -272 2409 -238
rect 2629 -272 2645 -238
rect 2851 -272 2867 -238
rect 3087 -272 3103 -238
rect 3309 -272 3325 -238
rect 3545 -272 3561 -238
rect -3815 -376 -3781 -314
rect 3781 -376 3815 -314
rect -3815 -410 -3719 -376
rect 3719 -410 3815 -376
<< viali >>
rect -3545 238 -3325 272
rect -3087 238 -2867 272
rect -2629 238 -2409 272
rect -2171 238 -1951 272
rect -1713 238 -1493 272
rect -1255 238 -1035 272
rect -797 238 -577 272
rect -339 238 -119 272
rect 119 238 339 272
rect 577 238 797 272
rect 1035 238 1255 272
rect 1493 238 1713 272
rect 1951 238 2171 272
rect 2409 238 2629 272
rect 2867 238 3087 272
rect 3325 238 3545 272
rect -3681 -188 -3647 188
rect -3223 -188 -3189 188
rect -2765 -188 -2731 188
rect -2307 -188 -2273 188
rect -1849 -188 -1815 188
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect 1815 -188 1849 188
rect 2273 -188 2307 188
rect 2731 -188 2765 188
rect 3189 -188 3223 188
rect 3647 -188 3681 188
rect -3545 -272 -3325 -238
rect -3087 -272 -2867 -238
rect -2629 -272 -2409 -238
rect -2171 -272 -1951 -238
rect -1713 -272 -1493 -238
rect -1255 -272 -1035 -238
rect -797 -272 -577 -238
rect -339 -272 -119 -238
rect 119 -272 339 -238
rect 577 -272 797 -238
rect 1035 -272 1255 -238
rect 1493 -272 1713 -238
rect 1951 -272 2171 -238
rect 2409 -272 2629 -238
rect 2867 -272 3087 -238
rect 3325 -272 3545 -238
<< metal1 >>
rect -3557 272 -3313 278
rect -3557 238 -3545 272
rect -3325 238 -3313 272
rect -3557 232 -3313 238
rect -3099 272 -2855 278
rect -3099 238 -3087 272
rect -2867 238 -2855 272
rect -3099 232 -2855 238
rect -2641 272 -2397 278
rect -2641 238 -2629 272
rect -2409 238 -2397 272
rect -2641 232 -2397 238
rect -2183 272 -1939 278
rect -2183 238 -2171 272
rect -1951 238 -1939 272
rect -2183 232 -1939 238
rect -1725 272 -1481 278
rect -1725 238 -1713 272
rect -1493 238 -1481 272
rect -1725 232 -1481 238
rect -1267 272 -1023 278
rect -1267 238 -1255 272
rect -1035 238 -1023 272
rect -1267 232 -1023 238
rect -809 272 -565 278
rect -809 238 -797 272
rect -577 238 -565 272
rect -809 232 -565 238
rect -351 272 -107 278
rect -351 238 -339 272
rect -119 238 -107 272
rect -351 232 -107 238
rect 107 272 351 278
rect 107 238 119 272
rect 339 238 351 272
rect 107 232 351 238
rect 565 272 809 278
rect 565 238 577 272
rect 797 238 809 272
rect 565 232 809 238
rect 1023 272 1267 278
rect 1023 238 1035 272
rect 1255 238 1267 272
rect 1023 232 1267 238
rect 1481 272 1725 278
rect 1481 238 1493 272
rect 1713 238 1725 272
rect 1481 232 1725 238
rect 1939 272 2183 278
rect 1939 238 1951 272
rect 2171 238 2183 272
rect 1939 232 2183 238
rect 2397 272 2641 278
rect 2397 238 2409 272
rect 2629 238 2641 272
rect 2397 232 2641 238
rect 2855 272 3099 278
rect 2855 238 2867 272
rect 3087 238 3099 272
rect 2855 232 3099 238
rect 3313 272 3557 278
rect 3313 238 3325 272
rect 3545 238 3557 272
rect 3313 232 3557 238
rect -3687 188 -3641 200
rect -3687 -188 -3681 188
rect -3647 -188 -3641 188
rect -3687 -200 -3641 -188
rect -3229 188 -3183 200
rect -3229 -188 -3223 188
rect -3189 -188 -3183 188
rect -3229 -200 -3183 -188
rect -2771 188 -2725 200
rect -2771 -188 -2765 188
rect -2731 -188 -2725 188
rect -2771 -200 -2725 -188
rect -2313 188 -2267 200
rect -2313 -188 -2307 188
rect -2273 -188 -2267 188
rect -2313 -200 -2267 -188
rect -1855 188 -1809 200
rect -1855 -188 -1849 188
rect -1815 -188 -1809 188
rect -1855 -200 -1809 -188
rect -1397 188 -1351 200
rect -1397 -188 -1391 188
rect -1357 -188 -1351 188
rect -1397 -200 -1351 -188
rect -939 188 -893 200
rect -939 -188 -933 188
rect -899 -188 -893 188
rect -939 -200 -893 -188
rect -481 188 -435 200
rect -481 -188 -475 188
rect -441 -188 -435 188
rect -481 -200 -435 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 435 188 481 200
rect 435 -188 441 188
rect 475 -188 481 188
rect 435 -200 481 -188
rect 893 188 939 200
rect 893 -188 899 188
rect 933 -188 939 188
rect 893 -200 939 -188
rect 1351 188 1397 200
rect 1351 -188 1357 188
rect 1391 -188 1397 188
rect 1351 -200 1397 -188
rect 1809 188 1855 200
rect 1809 -188 1815 188
rect 1849 -188 1855 188
rect 1809 -200 1855 -188
rect 2267 188 2313 200
rect 2267 -188 2273 188
rect 2307 -188 2313 188
rect 2267 -200 2313 -188
rect 2725 188 2771 200
rect 2725 -188 2731 188
rect 2765 -188 2771 188
rect 2725 -200 2771 -188
rect 3183 188 3229 200
rect 3183 -188 3189 188
rect 3223 -188 3229 188
rect 3183 -200 3229 -188
rect 3641 188 3687 200
rect 3641 -188 3647 188
rect 3681 -188 3687 188
rect 3641 -200 3687 -188
rect -3557 -238 -3313 -232
rect -3557 -272 -3545 -238
rect -3325 -272 -3313 -238
rect -3557 -278 -3313 -272
rect -3099 -238 -2855 -232
rect -3099 -272 -3087 -238
rect -2867 -272 -2855 -238
rect -3099 -278 -2855 -272
rect -2641 -238 -2397 -232
rect -2641 -272 -2629 -238
rect -2409 -272 -2397 -238
rect -2641 -278 -2397 -272
rect -2183 -238 -1939 -232
rect -2183 -272 -2171 -238
rect -1951 -272 -1939 -238
rect -2183 -278 -1939 -272
rect -1725 -238 -1481 -232
rect -1725 -272 -1713 -238
rect -1493 -272 -1481 -238
rect -1725 -278 -1481 -272
rect -1267 -238 -1023 -232
rect -1267 -272 -1255 -238
rect -1035 -272 -1023 -238
rect -1267 -278 -1023 -272
rect -809 -238 -565 -232
rect -809 -272 -797 -238
rect -577 -272 -565 -238
rect -809 -278 -565 -272
rect -351 -238 -107 -232
rect -351 -272 -339 -238
rect -119 -272 -107 -238
rect -351 -278 -107 -272
rect 107 -238 351 -232
rect 107 -272 119 -238
rect 339 -272 351 -238
rect 107 -278 351 -272
rect 565 -238 809 -232
rect 565 -272 577 -238
rect 797 -272 809 -238
rect 565 -278 809 -272
rect 1023 -238 1267 -232
rect 1023 -272 1035 -238
rect 1255 -272 1267 -238
rect 1023 -278 1267 -272
rect 1481 -238 1725 -232
rect 1481 -272 1493 -238
rect 1713 -272 1725 -238
rect 1481 -278 1725 -272
rect 1939 -238 2183 -232
rect 1939 -272 1951 -238
rect 2171 -272 2183 -238
rect 1939 -278 2183 -272
rect 2397 -238 2641 -232
rect 2397 -272 2409 -238
rect 2629 -272 2641 -238
rect 2397 -278 2641 -272
rect 2855 -238 3099 -232
rect 2855 -272 2867 -238
rect 3087 -272 3099 -238
rect 2855 -278 3099 -272
rect 3313 -238 3557 -232
rect 3313 -272 3325 -238
rect 3545 -272 3557 -238
rect 3313 -278 3557 -272
<< properties >>
string FIXED_BBOX -3798 -393 3798 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 16 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713232886
<< pwell >>
rect -3521 -810 3521 810
<< nmos >>
rect -3325 -600 -3125 600
rect -3067 -600 -2867 600
rect -2809 -600 -2609 600
rect -2551 -600 -2351 600
rect -2293 -600 -2093 600
rect -2035 -600 -1835 600
rect -1777 -600 -1577 600
rect -1519 -600 -1319 600
rect -1261 -600 -1061 600
rect -1003 -600 -803 600
rect -745 -600 -545 600
rect -487 -600 -287 600
rect -229 -600 -29 600
rect 29 -600 229 600
rect 287 -600 487 600
rect 545 -600 745 600
rect 803 -600 1003 600
rect 1061 -600 1261 600
rect 1319 -600 1519 600
rect 1577 -600 1777 600
rect 1835 -600 2035 600
rect 2093 -600 2293 600
rect 2351 -600 2551 600
rect 2609 -600 2809 600
rect 2867 -600 3067 600
rect 3125 -600 3325 600
<< ndiff >>
rect -3383 588 -3325 600
rect -3383 -588 -3371 588
rect -3337 -588 -3325 588
rect -3383 -600 -3325 -588
rect -3125 588 -3067 600
rect -3125 -588 -3113 588
rect -3079 -588 -3067 588
rect -3125 -600 -3067 -588
rect -2867 588 -2809 600
rect -2867 -588 -2855 588
rect -2821 -588 -2809 588
rect -2867 -600 -2809 -588
rect -2609 588 -2551 600
rect -2609 -588 -2597 588
rect -2563 -588 -2551 588
rect -2609 -600 -2551 -588
rect -2351 588 -2293 600
rect -2351 -588 -2339 588
rect -2305 -588 -2293 588
rect -2351 -600 -2293 -588
rect -2093 588 -2035 600
rect -2093 -588 -2081 588
rect -2047 -588 -2035 588
rect -2093 -600 -2035 -588
rect -1835 588 -1777 600
rect -1835 -588 -1823 588
rect -1789 -588 -1777 588
rect -1835 -600 -1777 -588
rect -1577 588 -1519 600
rect -1577 -588 -1565 588
rect -1531 -588 -1519 588
rect -1577 -600 -1519 -588
rect -1319 588 -1261 600
rect -1319 -588 -1307 588
rect -1273 -588 -1261 588
rect -1319 -600 -1261 -588
rect -1061 588 -1003 600
rect -1061 -588 -1049 588
rect -1015 -588 -1003 588
rect -1061 -600 -1003 -588
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -545 588 -487 600
rect -545 -588 -533 588
rect -499 -588 -487 588
rect -545 -600 -487 -588
rect -287 588 -229 600
rect -287 -588 -275 588
rect -241 -588 -229 588
rect -287 -600 -229 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 229 588 287 600
rect 229 -588 241 588
rect 275 -588 287 588
rect 229 -600 287 -588
rect 487 588 545 600
rect 487 -588 499 588
rect 533 -588 545 588
rect 487 -600 545 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
rect 1003 588 1061 600
rect 1003 -588 1015 588
rect 1049 -588 1061 588
rect 1003 -600 1061 -588
rect 1261 588 1319 600
rect 1261 -588 1273 588
rect 1307 -588 1319 588
rect 1261 -600 1319 -588
rect 1519 588 1577 600
rect 1519 -588 1531 588
rect 1565 -588 1577 588
rect 1519 -600 1577 -588
rect 1777 588 1835 600
rect 1777 -588 1789 588
rect 1823 -588 1835 588
rect 1777 -600 1835 -588
rect 2035 588 2093 600
rect 2035 -588 2047 588
rect 2081 -588 2093 588
rect 2035 -600 2093 -588
rect 2293 588 2351 600
rect 2293 -588 2305 588
rect 2339 -588 2351 588
rect 2293 -600 2351 -588
rect 2551 588 2609 600
rect 2551 -588 2563 588
rect 2597 -588 2609 588
rect 2551 -600 2609 -588
rect 2809 588 2867 600
rect 2809 -588 2821 588
rect 2855 -588 2867 588
rect 2809 -600 2867 -588
rect 3067 588 3125 600
rect 3067 -588 3079 588
rect 3113 -588 3125 588
rect 3067 -600 3125 -588
rect 3325 588 3383 600
rect 3325 -588 3337 588
rect 3371 -588 3383 588
rect 3325 -600 3383 -588
<< ndiffc >>
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
<< psubdiff >>
rect -3485 740 -3389 774
rect 3389 740 3485 774
rect -3485 678 -3451 740
rect 3451 678 3485 740
rect -3485 -740 -3451 -678
rect 3451 -740 3485 -678
rect -3485 -774 -3389 -740
rect 3389 -774 3485 -740
<< psubdiffcont >>
rect -3389 740 3389 774
rect -3485 -678 -3451 678
rect 3451 -678 3485 678
rect -3389 -774 3389 -740
<< poly >>
rect -3325 672 -3125 688
rect -3325 638 -3309 672
rect -3141 638 -3125 672
rect -3325 600 -3125 638
rect -3067 672 -2867 688
rect -3067 638 -3051 672
rect -2883 638 -2867 672
rect -3067 600 -2867 638
rect -2809 672 -2609 688
rect -2809 638 -2793 672
rect -2625 638 -2609 672
rect -2809 600 -2609 638
rect -2551 672 -2351 688
rect -2551 638 -2535 672
rect -2367 638 -2351 672
rect -2551 600 -2351 638
rect -2293 672 -2093 688
rect -2293 638 -2277 672
rect -2109 638 -2093 672
rect -2293 600 -2093 638
rect -2035 672 -1835 688
rect -2035 638 -2019 672
rect -1851 638 -1835 672
rect -2035 600 -1835 638
rect -1777 672 -1577 688
rect -1777 638 -1761 672
rect -1593 638 -1577 672
rect -1777 600 -1577 638
rect -1519 672 -1319 688
rect -1519 638 -1503 672
rect -1335 638 -1319 672
rect -1519 600 -1319 638
rect -1261 672 -1061 688
rect -1261 638 -1245 672
rect -1077 638 -1061 672
rect -1261 600 -1061 638
rect -1003 672 -803 688
rect -1003 638 -987 672
rect -819 638 -803 672
rect -1003 600 -803 638
rect -745 672 -545 688
rect -745 638 -729 672
rect -561 638 -545 672
rect -745 600 -545 638
rect -487 672 -287 688
rect -487 638 -471 672
rect -303 638 -287 672
rect -487 600 -287 638
rect -229 672 -29 688
rect -229 638 -213 672
rect -45 638 -29 672
rect -229 600 -29 638
rect 29 672 229 688
rect 29 638 45 672
rect 213 638 229 672
rect 29 600 229 638
rect 287 672 487 688
rect 287 638 303 672
rect 471 638 487 672
rect 287 600 487 638
rect 545 672 745 688
rect 545 638 561 672
rect 729 638 745 672
rect 545 600 745 638
rect 803 672 1003 688
rect 803 638 819 672
rect 987 638 1003 672
rect 803 600 1003 638
rect 1061 672 1261 688
rect 1061 638 1077 672
rect 1245 638 1261 672
rect 1061 600 1261 638
rect 1319 672 1519 688
rect 1319 638 1335 672
rect 1503 638 1519 672
rect 1319 600 1519 638
rect 1577 672 1777 688
rect 1577 638 1593 672
rect 1761 638 1777 672
rect 1577 600 1777 638
rect 1835 672 2035 688
rect 1835 638 1851 672
rect 2019 638 2035 672
rect 1835 600 2035 638
rect 2093 672 2293 688
rect 2093 638 2109 672
rect 2277 638 2293 672
rect 2093 600 2293 638
rect 2351 672 2551 688
rect 2351 638 2367 672
rect 2535 638 2551 672
rect 2351 600 2551 638
rect 2609 672 2809 688
rect 2609 638 2625 672
rect 2793 638 2809 672
rect 2609 600 2809 638
rect 2867 672 3067 688
rect 2867 638 2883 672
rect 3051 638 3067 672
rect 2867 600 3067 638
rect 3125 672 3325 688
rect 3125 638 3141 672
rect 3309 638 3325 672
rect 3125 600 3325 638
rect -3325 -638 -3125 -600
rect -3325 -672 -3309 -638
rect -3141 -672 -3125 -638
rect -3325 -688 -3125 -672
rect -3067 -638 -2867 -600
rect -3067 -672 -3051 -638
rect -2883 -672 -2867 -638
rect -3067 -688 -2867 -672
rect -2809 -638 -2609 -600
rect -2809 -672 -2793 -638
rect -2625 -672 -2609 -638
rect -2809 -688 -2609 -672
rect -2551 -638 -2351 -600
rect -2551 -672 -2535 -638
rect -2367 -672 -2351 -638
rect -2551 -688 -2351 -672
rect -2293 -638 -2093 -600
rect -2293 -672 -2277 -638
rect -2109 -672 -2093 -638
rect -2293 -688 -2093 -672
rect -2035 -638 -1835 -600
rect -2035 -672 -2019 -638
rect -1851 -672 -1835 -638
rect -2035 -688 -1835 -672
rect -1777 -638 -1577 -600
rect -1777 -672 -1761 -638
rect -1593 -672 -1577 -638
rect -1777 -688 -1577 -672
rect -1519 -638 -1319 -600
rect -1519 -672 -1503 -638
rect -1335 -672 -1319 -638
rect -1519 -688 -1319 -672
rect -1261 -638 -1061 -600
rect -1261 -672 -1245 -638
rect -1077 -672 -1061 -638
rect -1261 -688 -1061 -672
rect -1003 -638 -803 -600
rect -1003 -672 -987 -638
rect -819 -672 -803 -638
rect -1003 -688 -803 -672
rect -745 -638 -545 -600
rect -745 -672 -729 -638
rect -561 -672 -545 -638
rect -745 -688 -545 -672
rect -487 -638 -287 -600
rect -487 -672 -471 -638
rect -303 -672 -287 -638
rect -487 -688 -287 -672
rect -229 -638 -29 -600
rect -229 -672 -213 -638
rect -45 -672 -29 -638
rect -229 -688 -29 -672
rect 29 -638 229 -600
rect 29 -672 45 -638
rect 213 -672 229 -638
rect 29 -688 229 -672
rect 287 -638 487 -600
rect 287 -672 303 -638
rect 471 -672 487 -638
rect 287 -688 487 -672
rect 545 -638 745 -600
rect 545 -672 561 -638
rect 729 -672 745 -638
rect 545 -688 745 -672
rect 803 -638 1003 -600
rect 803 -672 819 -638
rect 987 -672 1003 -638
rect 803 -688 1003 -672
rect 1061 -638 1261 -600
rect 1061 -672 1077 -638
rect 1245 -672 1261 -638
rect 1061 -688 1261 -672
rect 1319 -638 1519 -600
rect 1319 -672 1335 -638
rect 1503 -672 1519 -638
rect 1319 -688 1519 -672
rect 1577 -638 1777 -600
rect 1577 -672 1593 -638
rect 1761 -672 1777 -638
rect 1577 -688 1777 -672
rect 1835 -638 2035 -600
rect 1835 -672 1851 -638
rect 2019 -672 2035 -638
rect 1835 -688 2035 -672
rect 2093 -638 2293 -600
rect 2093 -672 2109 -638
rect 2277 -672 2293 -638
rect 2093 -688 2293 -672
rect 2351 -638 2551 -600
rect 2351 -672 2367 -638
rect 2535 -672 2551 -638
rect 2351 -688 2551 -672
rect 2609 -638 2809 -600
rect 2609 -672 2625 -638
rect 2793 -672 2809 -638
rect 2609 -688 2809 -672
rect 2867 -638 3067 -600
rect 2867 -672 2883 -638
rect 3051 -672 3067 -638
rect 2867 -688 3067 -672
rect 3125 -638 3325 -600
rect 3125 -672 3141 -638
rect 3309 -672 3325 -638
rect 3125 -688 3325 -672
<< polycont >>
rect -3309 638 -3141 672
rect -3051 638 -2883 672
rect -2793 638 -2625 672
rect -2535 638 -2367 672
rect -2277 638 -2109 672
rect -2019 638 -1851 672
rect -1761 638 -1593 672
rect -1503 638 -1335 672
rect -1245 638 -1077 672
rect -987 638 -819 672
rect -729 638 -561 672
rect -471 638 -303 672
rect -213 638 -45 672
rect 45 638 213 672
rect 303 638 471 672
rect 561 638 729 672
rect 819 638 987 672
rect 1077 638 1245 672
rect 1335 638 1503 672
rect 1593 638 1761 672
rect 1851 638 2019 672
rect 2109 638 2277 672
rect 2367 638 2535 672
rect 2625 638 2793 672
rect 2883 638 3051 672
rect 3141 638 3309 672
rect -3309 -672 -3141 -638
rect -3051 -672 -2883 -638
rect -2793 -672 -2625 -638
rect -2535 -672 -2367 -638
rect -2277 -672 -2109 -638
rect -2019 -672 -1851 -638
rect -1761 -672 -1593 -638
rect -1503 -672 -1335 -638
rect -1245 -672 -1077 -638
rect -987 -672 -819 -638
rect -729 -672 -561 -638
rect -471 -672 -303 -638
rect -213 -672 -45 -638
rect 45 -672 213 -638
rect 303 -672 471 -638
rect 561 -672 729 -638
rect 819 -672 987 -638
rect 1077 -672 1245 -638
rect 1335 -672 1503 -638
rect 1593 -672 1761 -638
rect 1851 -672 2019 -638
rect 2109 -672 2277 -638
rect 2367 -672 2535 -638
rect 2625 -672 2793 -638
rect 2883 -672 3051 -638
rect 3141 -672 3309 -638
<< locali >>
rect -3485 740 -3389 774
rect 3389 740 3485 774
rect -3485 678 -3451 740
rect 3451 678 3485 740
rect -3325 638 -3309 672
rect -3141 638 -3125 672
rect -3067 638 -3051 672
rect -2883 638 -2867 672
rect -2809 638 -2793 672
rect -2625 638 -2609 672
rect -2551 638 -2535 672
rect -2367 638 -2351 672
rect -2293 638 -2277 672
rect -2109 638 -2093 672
rect -2035 638 -2019 672
rect -1851 638 -1835 672
rect -1777 638 -1761 672
rect -1593 638 -1577 672
rect -1519 638 -1503 672
rect -1335 638 -1319 672
rect -1261 638 -1245 672
rect -1077 638 -1061 672
rect -1003 638 -987 672
rect -819 638 -803 672
rect -745 638 -729 672
rect -561 638 -545 672
rect -487 638 -471 672
rect -303 638 -287 672
rect -229 638 -213 672
rect -45 638 -29 672
rect 29 638 45 672
rect 213 638 229 672
rect 287 638 303 672
rect 471 638 487 672
rect 545 638 561 672
rect 729 638 745 672
rect 803 638 819 672
rect 987 638 1003 672
rect 1061 638 1077 672
rect 1245 638 1261 672
rect 1319 638 1335 672
rect 1503 638 1519 672
rect 1577 638 1593 672
rect 1761 638 1777 672
rect 1835 638 1851 672
rect 2019 638 2035 672
rect 2093 638 2109 672
rect 2277 638 2293 672
rect 2351 638 2367 672
rect 2535 638 2551 672
rect 2609 638 2625 672
rect 2793 638 2809 672
rect 2867 638 2883 672
rect 3051 638 3067 672
rect 3125 638 3141 672
rect 3309 638 3325 672
rect -3371 588 -3337 604
rect -3371 -604 -3337 -588
rect -3113 588 -3079 604
rect -3113 -604 -3079 -588
rect -2855 588 -2821 604
rect -2855 -604 -2821 -588
rect -2597 588 -2563 604
rect -2597 -604 -2563 -588
rect -2339 588 -2305 604
rect -2339 -604 -2305 -588
rect -2081 588 -2047 604
rect -2081 -604 -2047 -588
rect -1823 588 -1789 604
rect -1823 -604 -1789 -588
rect -1565 588 -1531 604
rect -1565 -604 -1531 -588
rect -1307 588 -1273 604
rect -1307 -604 -1273 -588
rect -1049 588 -1015 604
rect -1049 -604 -1015 -588
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -533 588 -499 604
rect -533 -604 -499 -588
rect -275 588 -241 604
rect -275 -604 -241 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 241 588 275 604
rect 241 -604 275 -588
rect 499 588 533 604
rect 499 -604 533 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect 1015 588 1049 604
rect 1015 -604 1049 -588
rect 1273 588 1307 604
rect 1273 -604 1307 -588
rect 1531 588 1565 604
rect 1531 -604 1565 -588
rect 1789 588 1823 604
rect 1789 -604 1823 -588
rect 2047 588 2081 604
rect 2047 -604 2081 -588
rect 2305 588 2339 604
rect 2305 -604 2339 -588
rect 2563 588 2597 604
rect 2563 -604 2597 -588
rect 2821 588 2855 604
rect 2821 -604 2855 -588
rect 3079 588 3113 604
rect 3079 -604 3113 -588
rect 3337 588 3371 604
rect 3337 -604 3371 -588
rect -3325 -672 -3309 -638
rect -3141 -672 -3125 -638
rect -3067 -672 -3051 -638
rect -2883 -672 -2867 -638
rect -2809 -672 -2793 -638
rect -2625 -672 -2609 -638
rect -2551 -672 -2535 -638
rect -2367 -672 -2351 -638
rect -2293 -672 -2277 -638
rect -2109 -672 -2093 -638
rect -2035 -672 -2019 -638
rect -1851 -672 -1835 -638
rect -1777 -672 -1761 -638
rect -1593 -672 -1577 -638
rect -1519 -672 -1503 -638
rect -1335 -672 -1319 -638
rect -1261 -672 -1245 -638
rect -1077 -672 -1061 -638
rect -1003 -672 -987 -638
rect -819 -672 -803 -638
rect -745 -672 -729 -638
rect -561 -672 -545 -638
rect -487 -672 -471 -638
rect -303 -672 -287 -638
rect -229 -672 -213 -638
rect -45 -672 -29 -638
rect 29 -672 45 -638
rect 213 -672 229 -638
rect 287 -672 303 -638
rect 471 -672 487 -638
rect 545 -672 561 -638
rect 729 -672 745 -638
rect 803 -672 819 -638
rect 987 -672 1003 -638
rect 1061 -672 1077 -638
rect 1245 -672 1261 -638
rect 1319 -672 1335 -638
rect 1503 -672 1519 -638
rect 1577 -672 1593 -638
rect 1761 -672 1777 -638
rect 1835 -672 1851 -638
rect 2019 -672 2035 -638
rect 2093 -672 2109 -638
rect 2277 -672 2293 -638
rect 2351 -672 2367 -638
rect 2535 -672 2551 -638
rect 2609 -672 2625 -638
rect 2793 -672 2809 -638
rect 2867 -672 2883 -638
rect 3051 -672 3067 -638
rect 3125 -672 3141 -638
rect 3309 -672 3325 -638
rect -3485 -740 -3451 -678
rect 3451 -740 3485 -678
rect -3485 -774 -3389 -740
rect 3389 -774 3485 -740
<< viali >>
rect -3309 638 -3141 672
rect -3051 638 -2883 672
rect -2793 638 -2625 672
rect -2535 638 -2367 672
rect -2277 638 -2109 672
rect -2019 638 -1851 672
rect -1761 638 -1593 672
rect -1503 638 -1335 672
rect -1245 638 -1077 672
rect -987 638 -819 672
rect -729 638 -561 672
rect -471 638 -303 672
rect -213 638 -45 672
rect 45 638 213 672
rect 303 638 471 672
rect 561 638 729 672
rect 819 638 987 672
rect 1077 638 1245 672
rect 1335 638 1503 672
rect 1593 638 1761 672
rect 1851 638 2019 672
rect 2109 638 2277 672
rect 2367 638 2535 672
rect 2625 638 2793 672
rect 2883 638 3051 672
rect 3141 638 3309 672
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
rect -3309 -672 -3141 -638
rect -3051 -672 -2883 -638
rect -2793 -672 -2625 -638
rect -2535 -672 -2367 -638
rect -2277 -672 -2109 -638
rect -2019 -672 -1851 -638
rect -1761 -672 -1593 -638
rect -1503 -672 -1335 -638
rect -1245 -672 -1077 -638
rect -987 -672 -819 -638
rect -729 -672 -561 -638
rect -471 -672 -303 -638
rect -213 -672 -45 -638
rect 45 -672 213 -638
rect 303 -672 471 -638
rect 561 -672 729 -638
rect 819 -672 987 -638
rect 1077 -672 1245 -638
rect 1335 -672 1503 -638
rect 1593 -672 1761 -638
rect 1851 -672 2019 -638
rect 2109 -672 2277 -638
rect 2367 -672 2535 -638
rect 2625 -672 2793 -638
rect 2883 -672 3051 -638
rect 3141 -672 3309 -638
<< metal1 >>
rect -3321 672 -3129 678
rect -3321 638 -3309 672
rect -3141 638 -3129 672
rect -3321 632 -3129 638
rect -3063 672 -2871 678
rect -3063 638 -3051 672
rect -2883 638 -2871 672
rect -3063 632 -2871 638
rect -2805 672 -2613 678
rect -2805 638 -2793 672
rect -2625 638 -2613 672
rect -2805 632 -2613 638
rect -2547 672 -2355 678
rect -2547 638 -2535 672
rect -2367 638 -2355 672
rect -2547 632 -2355 638
rect -2289 672 -2097 678
rect -2289 638 -2277 672
rect -2109 638 -2097 672
rect -2289 632 -2097 638
rect -2031 672 -1839 678
rect -2031 638 -2019 672
rect -1851 638 -1839 672
rect -2031 632 -1839 638
rect -1773 672 -1581 678
rect -1773 638 -1761 672
rect -1593 638 -1581 672
rect -1773 632 -1581 638
rect -1515 672 -1323 678
rect -1515 638 -1503 672
rect -1335 638 -1323 672
rect -1515 632 -1323 638
rect -1257 672 -1065 678
rect -1257 638 -1245 672
rect -1077 638 -1065 672
rect -1257 632 -1065 638
rect -999 672 -807 678
rect -999 638 -987 672
rect -819 638 -807 672
rect -999 632 -807 638
rect -741 672 -549 678
rect -741 638 -729 672
rect -561 638 -549 672
rect -741 632 -549 638
rect -483 672 -291 678
rect -483 638 -471 672
rect -303 638 -291 672
rect -483 632 -291 638
rect -225 672 -33 678
rect -225 638 -213 672
rect -45 638 -33 672
rect -225 632 -33 638
rect 33 672 225 678
rect 33 638 45 672
rect 213 638 225 672
rect 33 632 225 638
rect 291 672 483 678
rect 291 638 303 672
rect 471 638 483 672
rect 291 632 483 638
rect 549 672 741 678
rect 549 638 561 672
rect 729 638 741 672
rect 549 632 741 638
rect 807 672 999 678
rect 807 638 819 672
rect 987 638 999 672
rect 807 632 999 638
rect 1065 672 1257 678
rect 1065 638 1077 672
rect 1245 638 1257 672
rect 1065 632 1257 638
rect 1323 672 1515 678
rect 1323 638 1335 672
rect 1503 638 1515 672
rect 1323 632 1515 638
rect 1581 672 1773 678
rect 1581 638 1593 672
rect 1761 638 1773 672
rect 1581 632 1773 638
rect 1839 672 2031 678
rect 1839 638 1851 672
rect 2019 638 2031 672
rect 1839 632 2031 638
rect 2097 672 2289 678
rect 2097 638 2109 672
rect 2277 638 2289 672
rect 2097 632 2289 638
rect 2355 672 2547 678
rect 2355 638 2367 672
rect 2535 638 2547 672
rect 2355 632 2547 638
rect 2613 672 2805 678
rect 2613 638 2625 672
rect 2793 638 2805 672
rect 2613 632 2805 638
rect 2871 672 3063 678
rect 2871 638 2883 672
rect 3051 638 3063 672
rect 2871 632 3063 638
rect 3129 672 3321 678
rect 3129 638 3141 672
rect 3309 638 3321 672
rect 3129 632 3321 638
rect -3377 588 -3331 600
rect -3377 -588 -3371 588
rect -3337 -588 -3331 588
rect -3377 -600 -3331 -588
rect -3119 588 -3073 600
rect -3119 -588 -3113 588
rect -3079 -588 -3073 588
rect -3119 -600 -3073 -588
rect -2861 588 -2815 600
rect -2861 -588 -2855 588
rect -2821 -588 -2815 588
rect -2861 -600 -2815 -588
rect -2603 588 -2557 600
rect -2603 -588 -2597 588
rect -2563 -588 -2557 588
rect -2603 -600 -2557 -588
rect -2345 588 -2299 600
rect -2345 -588 -2339 588
rect -2305 -588 -2299 588
rect -2345 -600 -2299 -588
rect -2087 588 -2041 600
rect -2087 -588 -2081 588
rect -2047 -588 -2041 588
rect -2087 -600 -2041 -588
rect -1829 588 -1783 600
rect -1829 -588 -1823 588
rect -1789 -588 -1783 588
rect -1829 -600 -1783 -588
rect -1571 588 -1525 600
rect -1571 -588 -1565 588
rect -1531 -588 -1525 588
rect -1571 -600 -1525 -588
rect -1313 588 -1267 600
rect -1313 -588 -1307 588
rect -1273 -588 -1267 588
rect -1313 -600 -1267 -588
rect -1055 588 -1009 600
rect -1055 -588 -1049 588
rect -1015 -588 -1009 588
rect -1055 -600 -1009 -588
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -539 588 -493 600
rect -539 -588 -533 588
rect -499 -588 -493 588
rect -539 -600 -493 -588
rect -281 588 -235 600
rect -281 -588 -275 588
rect -241 -588 -235 588
rect -281 -600 -235 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 235 588 281 600
rect 235 -588 241 588
rect 275 -588 281 588
rect 235 -600 281 -588
rect 493 588 539 600
rect 493 -588 499 588
rect 533 -588 539 588
rect 493 -600 539 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect 1009 588 1055 600
rect 1009 -588 1015 588
rect 1049 -588 1055 588
rect 1009 -600 1055 -588
rect 1267 588 1313 600
rect 1267 -588 1273 588
rect 1307 -588 1313 588
rect 1267 -600 1313 -588
rect 1525 588 1571 600
rect 1525 -588 1531 588
rect 1565 -588 1571 588
rect 1525 -600 1571 -588
rect 1783 588 1829 600
rect 1783 -588 1789 588
rect 1823 -588 1829 588
rect 1783 -600 1829 -588
rect 2041 588 2087 600
rect 2041 -588 2047 588
rect 2081 -588 2087 588
rect 2041 -600 2087 -588
rect 2299 588 2345 600
rect 2299 -588 2305 588
rect 2339 -588 2345 588
rect 2299 -600 2345 -588
rect 2557 588 2603 600
rect 2557 -588 2563 588
rect 2597 -588 2603 588
rect 2557 -600 2603 -588
rect 2815 588 2861 600
rect 2815 -588 2821 588
rect 2855 -588 2861 588
rect 2815 -600 2861 -588
rect 3073 588 3119 600
rect 3073 -588 3079 588
rect 3113 -588 3119 588
rect 3073 -600 3119 -588
rect 3331 588 3377 600
rect 3331 -588 3337 588
rect 3371 -588 3377 588
rect 3331 -600 3377 -588
rect -3321 -638 -3129 -632
rect -3321 -672 -3309 -638
rect -3141 -672 -3129 -638
rect -3321 -678 -3129 -672
rect -3063 -638 -2871 -632
rect -3063 -672 -3051 -638
rect -2883 -672 -2871 -638
rect -3063 -678 -2871 -672
rect -2805 -638 -2613 -632
rect -2805 -672 -2793 -638
rect -2625 -672 -2613 -638
rect -2805 -678 -2613 -672
rect -2547 -638 -2355 -632
rect -2547 -672 -2535 -638
rect -2367 -672 -2355 -638
rect -2547 -678 -2355 -672
rect -2289 -638 -2097 -632
rect -2289 -672 -2277 -638
rect -2109 -672 -2097 -638
rect -2289 -678 -2097 -672
rect -2031 -638 -1839 -632
rect -2031 -672 -2019 -638
rect -1851 -672 -1839 -638
rect -2031 -678 -1839 -672
rect -1773 -638 -1581 -632
rect -1773 -672 -1761 -638
rect -1593 -672 -1581 -638
rect -1773 -678 -1581 -672
rect -1515 -638 -1323 -632
rect -1515 -672 -1503 -638
rect -1335 -672 -1323 -638
rect -1515 -678 -1323 -672
rect -1257 -638 -1065 -632
rect -1257 -672 -1245 -638
rect -1077 -672 -1065 -638
rect -1257 -678 -1065 -672
rect -999 -638 -807 -632
rect -999 -672 -987 -638
rect -819 -672 -807 -638
rect -999 -678 -807 -672
rect -741 -638 -549 -632
rect -741 -672 -729 -638
rect -561 -672 -549 -638
rect -741 -678 -549 -672
rect -483 -638 -291 -632
rect -483 -672 -471 -638
rect -303 -672 -291 -638
rect -483 -678 -291 -672
rect -225 -638 -33 -632
rect -225 -672 -213 -638
rect -45 -672 -33 -638
rect -225 -678 -33 -672
rect 33 -638 225 -632
rect 33 -672 45 -638
rect 213 -672 225 -638
rect 33 -678 225 -672
rect 291 -638 483 -632
rect 291 -672 303 -638
rect 471 -672 483 -638
rect 291 -678 483 -672
rect 549 -638 741 -632
rect 549 -672 561 -638
rect 729 -672 741 -638
rect 549 -678 741 -672
rect 807 -638 999 -632
rect 807 -672 819 -638
rect 987 -672 999 -638
rect 807 -678 999 -672
rect 1065 -638 1257 -632
rect 1065 -672 1077 -638
rect 1245 -672 1257 -638
rect 1065 -678 1257 -672
rect 1323 -638 1515 -632
rect 1323 -672 1335 -638
rect 1503 -672 1515 -638
rect 1323 -678 1515 -672
rect 1581 -638 1773 -632
rect 1581 -672 1593 -638
rect 1761 -672 1773 -638
rect 1581 -678 1773 -672
rect 1839 -638 2031 -632
rect 1839 -672 1851 -638
rect 2019 -672 2031 -638
rect 1839 -678 2031 -672
rect 2097 -638 2289 -632
rect 2097 -672 2109 -638
rect 2277 -672 2289 -638
rect 2097 -678 2289 -672
rect 2355 -638 2547 -632
rect 2355 -672 2367 -638
rect 2535 -672 2547 -638
rect 2355 -678 2547 -672
rect 2613 -638 2805 -632
rect 2613 -672 2625 -638
rect 2793 -672 2805 -638
rect 2613 -678 2805 -672
rect 2871 -638 3063 -632
rect 2871 -672 2883 -638
rect 3051 -672 3063 -638
rect 2871 -678 3063 -672
rect 3129 -638 3321 -632
rect 3129 -672 3141 -638
rect 3309 -672 3321 -638
rect 3129 -678 3321 -672
<< properties >>
string FIXED_BBOX -3468 -757 3468 757
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6 l 1 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

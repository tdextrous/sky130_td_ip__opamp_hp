magic
tech sky130A
magscale 1 2
timestamp 1713393625
<< nwell >>
rect -5389 -1497 5389 1497
<< mvpmos >>
rect -5131 -1200 -4931 1200
rect -4873 -1200 -4673 1200
rect -4615 -1200 -4415 1200
rect -4357 -1200 -4157 1200
rect -4099 -1200 -3899 1200
rect -3841 -1200 -3641 1200
rect -3583 -1200 -3383 1200
rect -3325 -1200 -3125 1200
rect -3067 -1200 -2867 1200
rect -2809 -1200 -2609 1200
rect -2551 -1200 -2351 1200
rect -2293 -1200 -2093 1200
rect -2035 -1200 -1835 1200
rect -1777 -1200 -1577 1200
rect -1519 -1200 -1319 1200
rect -1261 -1200 -1061 1200
rect -1003 -1200 -803 1200
rect -745 -1200 -545 1200
rect -487 -1200 -287 1200
rect -229 -1200 -29 1200
rect 29 -1200 229 1200
rect 287 -1200 487 1200
rect 545 -1200 745 1200
rect 803 -1200 1003 1200
rect 1061 -1200 1261 1200
rect 1319 -1200 1519 1200
rect 1577 -1200 1777 1200
rect 1835 -1200 2035 1200
rect 2093 -1200 2293 1200
rect 2351 -1200 2551 1200
rect 2609 -1200 2809 1200
rect 2867 -1200 3067 1200
rect 3125 -1200 3325 1200
rect 3383 -1200 3583 1200
rect 3641 -1200 3841 1200
rect 3899 -1200 4099 1200
rect 4157 -1200 4357 1200
rect 4415 -1200 4615 1200
rect 4673 -1200 4873 1200
rect 4931 -1200 5131 1200
<< mvpdiff >>
rect -5189 1188 -5131 1200
rect -5189 -1188 -5177 1188
rect -5143 -1188 -5131 1188
rect -5189 -1200 -5131 -1188
rect -4931 1188 -4873 1200
rect -4931 -1188 -4919 1188
rect -4885 -1188 -4873 1188
rect -4931 -1200 -4873 -1188
rect -4673 1188 -4615 1200
rect -4673 -1188 -4661 1188
rect -4627 -1188 -4615 1188
rect -4673 -1200 -4615 -1188
rect -4415 1188 -4357 1200
rect -4415 -1188 -4403 1188
rect -4369 -1188 -4357 1188
rect -4415 -1200 -4357 -1188
rect -4157 1188 -4099 1200
rect -4157 -1188 -4145 1188
rect -4111 -1188 -4099 1188
rect -4157 -1200 -4099 -1188
rect -3899 1188 -3841 1200
rect -3899 -1188 -3887 1188
rect -3853 -1188 -3841 1188
rect -3899 -1200 -3841 -1188
rect -3641 1188 -3583 1200
rect -3641 -1188 -3629 1188
rect -3595 -1188 -3583 1188
rect -3641 -1200 -3583 -1188
rect -3383 1188 -3325 1200
rect -3383 -1188 -3371 1188
rect -3337 -1188 -3325 1188
rect -3383 -1200 -3325 -1188
rect -3125 1188 -3067 1200
rect -3125 -1188 -3113 1188
rect -3079 -1188 -3067 1188
rect -3125 -1200 -3067 -1188
rect -2867 1188 -2809 1200
rect -2867 -1188 -2855 1188
rect -2821 -1188 -2809 1188
rect -2867 -1200 -2809 -1188
rect -2609 1188 -2551 1200
rect -2609 -1188 -2597 1188
rect -2563 -1188 -2551 1188
rect -2609 -1200 -2551 -1188
rect -2351 1188 -2293 1200
rect -2351 -1188 -2339 1188
rect -2305 -1188 -2293 1188
rect -2351 -1200 -2293 -1188
rect -2093 1188 -2035 1200
rect -2093 -1188 -2081 1188
rect -2047 -1188 -2035 1188
rect -2093 -1200 -2035 -1188
rect -1835 1188 -1777 1200
rect -1835 -1188 -1823 1188
rect -1789 -1188 -1777 1188
rect -1835 -1200 -1777 -1188
rect -1577 1188 -1519 1200
rect -1577 -1188 -1565 1188
rect -1531 -1188 -1519 1188
rect -1577 -1200 -1519 -1188
rect -1319 1188 -1261 1200
rect -1319 -1188 -1307 1188
rect -1273 -1188 -1261 1188
rect -1319 -1200 -1261 -1188
rect -1061 1188 -1003 1200
rect -1061 -1188 -1049 1188
rect -1015 -1188 -1003 1188
rect -1061 -1200 -1003 -1188
rect -803 1188 -745 1200
rect -803 -1188 -791 1188
rect -757 -1188 -745 1188
rect -803 -1200 -745 -1188
rect -545 1188 -487 1200
rect -545 -1188 -533 1188
rect -499 -1188 -487 1188
rect -545 -1200 -487 -1188
rect -287 1188 -229 1200
rect -287 -1188 -275 1188
rect -241 -1188 -229 1188
rect -287 -1200 -229 -1188
rect -29 1188 29 1200
rect -29 -1188 -17 1188
rect 17 -1188 29 1188
rect -29 -1200 29 -1188
rect 229 1188 287 1200
rect 229 -1188 241 1188
rect 275 -1188 287 1188
rect 229 -1200 287 -1188
rect 487 1188 545 1200
rect 487 -1188 499 1188
rect 533 -1188 545 1188
rect 487 -1200 545 -1188
rect 745 1188 803 1200
rect 745 -1188 757 1188
rect 791 -1188 803 1188
rect 745 -1200 803 -1188
rect 1003 1188 1061 1200
rect 1003 -1188 1015 1188
rect 1049 -1188 1061 1188
rect 1003 -1200 1061 -1188
rect 1261 1188 1319 1200
rect 1261 -1188 1273 1188
rect 1307 -1188 1319 1188
rect 1261 -1200 1319 -1188
rect 1519 1188 1577 1200
rect 1519 -1188 1531 1188
rect 1565 -1188 1577 1188
rect 1519 -1200 1577 -1188
rect 1777 1188 1835 1200
rect 1777 -1188 1789 1188
rect 1823 -1188 1835 1188
rect 1777 -1200 1835 -1188
rect 2035 1188 2093 1200
rect 2035 -1188 2047 1188
rect 2081 -1188 2093 1188
rect 2035 -1200 2093 -1188
rect 2293 1188 2351 1200
rect 2293 -1188 2305 1188
rect 2339 -1188 2351 1188
rect 2293 -1200 2351 -1188
rect 2551 1188 2609 1200
rect 2551 -1188 2563 1188
rect 2597 -1188 2609 1188
rect 2551 -1200 2609 -1188
rect 2809 1188 2867 1200
rect 2809 -1188 2821 1188
rect 2855 -1188 2867 1188
rect 2809 -1200 2867 -1188
rect 3067 1188 3125 1200
rect 3067 -1188 3079 1188
rect 3113 -1188 3125 1188
rect 3067 -1200 3125 -1188
rect 3325 1188 3383 1200
rect 3325 -1188 3337 1188
rect 3371 -1188 3383 1188
rect 3325 -1200 3383 -1188
rect 3583 1188 3641 1200
rect 3583 -1188 3595 1188
rect 3629 -1188 3641 1188
rect 3583 -1200 3641 -1188
rect 3841 1188 3899 1200
rect 3841 -1188 3853 1188
rect 3887 -1188 3899 1188
rect 3841 -1200 3899 -1188
rect 4099 1188 4157 1200
rect 4099 -1188 4111 1188
rect 4145 -1188 4157 1188
rect 4099 -1200 4157 -1188
rect 4357 1188 4415 1200
rect 4357 -1188 4369 1188
rect 4403 -1188 4415 1188
rect 4357 -1200 4415 -1188
rect 4615 1188 4673 1200
rect 4615 -1188 4627 1188
rect 4661 -1188 4673 1188
rect 4615 -1200 4673 -1188
rect 4873 1188 4931 1200
rect 4873 -1188 4885 1188
rect 4919 -1188 4931 1188
rect 4873 -1200 4931 -1188
rect 5131 1188 5189 1200
rect 5131 -1188 5143 1188
rect 5177 -1188 5189 1188
rect 5131 -1200 5189 -1188
<< mvpdiffc >>
rect -5177 -1188 -5143 1188
rect -4919 -1188 -4885 1188
rect -4661 -1188 -4627 1188
rect -4403 -1188 -4369 1188
rect -4145 -1188 -4111 1188
rect -3887 -1188 -3853 1188
rect -3629 -1188 -3595 1188
rect -3371 -1188 -3337 1188
rect -3113 -1188 -3079 1188
rect -2855 -1188 -2821 1188
rect -2597 -1188 -2563 1188
rect -2339 -1188 -2305 1188
rect -2081 -1188 -2047 1188
rect -1823 -1188 -1789 1188
rect -1565 -1188 -1531 1188
rect -1307 -1188 -1273 1188
rect -1049 -1188 -1015 1188
rect -791 -1188 -757 1188
rect -533 -1188 -499 1188
rect -275 -1188 -241 1188
rect -17 -1188 17 1188
rect 241 -1188 275 1188
rect 499 -1188 533 1188
rect 757 -1188 791 1188
rect 1015 -1188 1049 1188
rect 1273 -1188 1307 1188
rect 1531 -1188 1565 1188
rect 1789 -1188 1823 1188
rect 2047 -1188 2081 1188
rect 2305 -1188 2339 1188
rect 2563 -1188 2597 1188
rect 2821 -1188 2855 1188
rect 3079 -1188 3113 1188
rect 3337 -1188 3371 1188
rect 3595 -1188 3629 1188
rect 3853 -1188 3887 1188
rect 4111 -1188 4145 1188
rect 4369 -1188 4403 1188
rect 4627 -1188 4661 1188
rect 4885 -1188 4919 1188
rect 5143 -1188 5177 1188
<< mvnsubdiff >>
rect -5323 1419 5323 1431
rect -5323 1385 -5215 1419
rect 5215 1385 5323 1419
rect -5323 1373 5323 1385
rect -5323 1323 -5265 1373
rect -5323 -1323 -5311 1323
rect -5277 -1323 -5265 1323
rect 5265 1323 5323 1373
rect -5323 -1373 -5265 -1323
rect 5265 -1323 5277 1323
rect 5311 -1323 5323 1323
rect 5265 -1373 5323 -1323
rect -5323 -1385 5323 -1373
rect -5323 -1419 -5215 -1385
rect 5215 -1419 5323 -1385
rect -5323 -1431 5323 -1419
<< mvnsubdiffcont >>
rect -5215 1385 5215 1419
rect -5311 -1323 -5277 1323
rect 5277 -1323 5311 1323
rect -5215 -1419 5215 -1385
<< poly >>
rect -5097 1281 -4965 1297
rect -5097 1264 -5081 1281
rect -5131 1247 -5081 1264
rect -4981 1264 -4965 1281
rect -4839 1281 -4707 1297
rect -4839 1264 -4823 1281
rect -4981 1247 -4931 1264
rect -5131 1200 -4931 1247
rect -4873 1247 -4823 1264
rect -4723 1264 -4707 1281
rect -4581 1281 -4449 1297
rect -4581 1264 -4565 1281
rect -4723 1247 -4673 1264
rect -4873 1200 -4673 1247
rect -4615 1247 -4565 1264
rect -4465 1264 -4449 1281
rect -4323 1281 -4191 1297
rect -4323 1264 -4307 1281
rect -4465 1247 -4415 1264
rect -4615 1200 -4415 1247
rect -4357 1247 -4307 1264
rect -4207 1264 -4191 1281
rect -4065 1281 -3933 1297
rect -4065 1264 -4049 1281
rect -4207 1247 -4157 1264
rect -4357 1200 -4157 1247
rect -4099 1247 -4049 1264
rect -3949 1264 -3933 1281
rect -3807 1281 -3675 1297
rect -3807 1264 -3791 1281
rect -3949 1247 -3899 1264
rect -4099 1200 -3899 1247
rect -3841 1247 -3791 1264
rect -3691 1264 -3675 1281
rect -3549 1281 -3417 1297
rect -3549 1264 -3533 1281
rect -3691 1247 -3641 1264
rect -3841 1200 -3641 1247
rect -3583 1247 -3533 1264
rect -3433 1264 -3417 1281
rect -3291 1281 -3159 1297
rect -3291 1264 -3275 1281
rect -3433 1247 -3383 1264
rect -3583 1200 -3383 1247
rect -3325 1247 -3275 1264
rect -3175 1264 -3159 1281
rect -3033 1281 -2901 1297
rect -3033 1264 -3017 1281
rect -3175 1247 -3125 1264
rect -3325 1200 -3125 1247
rect -3067 1247 -3017 1264
rect -2917 1264 -2901 1281
rect -2775 1281 -2643 1297
rect -2775 1264 -2759 1281
rect -2917 1247 -2867 1264
rect -3067 1200 -2867 1247
rect -2809 1247 -2759 1264
rect -2659 1264 -2643 1281
rect -2517 1281 -2385 1297
rect -2517 1264 -2501 1281
rect -2659 1247 -2609 1264
rect -2809 1200 -2609 1247
rect -2551 1247 -2501 1264
rect -2401 1264 -2385 1281
rect -2259 1281 -2127 1297
rect -2259 1264 -2243 1281
rect -2401 1247 -2351 1264
rect -2551 1200 -2351 1247
rect -2293 1247 -2243 1264
rect -2143 1264 -2127 1281
rect -2001 1281 -1869 1297
rect -2001 1264 -1985 1281
rect -2143 1247 -2093 1264
rect -2293 1200 -2093 1247
rect -2035 1247 -1985 1264
rect -1885 1264 -1869 1281
rect -1743 1281 -1611 1297
rect -1743 1264 -1727 1281
rect -1885 1247 -1835 1264
rect -2035 1200 -1835 1247
rect -1777 1247 -1727 1264
rect -1627 1264 -1611 1281
rect -1485 1281 -1353 1297
rect -1485 1264 -1469 1281
rect -1627 1247 -1577 1264
rect -1777 1200 -1577 1247
rect -1519 1247 -1469 1264
rect -1369 1264 -1353 1281
rect -1227 1281 -1095 1297
rect -1227 1264 -1211 1281
rect -1369 1247 -1319 1264
rect -1519 1200 -1319 1247
rect -1261 1247 -1211 1264
rect -1111 1264 -1095 1281
rect -969 1281 -837 1297
rect -969 1264 -953 1281
rect -1111 1247 -1061 1264
rect -1261 1200 -1061 1247
rect -1003 1247 -953 1264
rect -853 1264 -837 1281
rect -711 1281 -579 1297
rect -711 1264 -695 1281
rect -853 1247 -803 1264
rect -1003 1200 -803 1247
rect -745 1247 -695 1264
rect -595 1264 -579 1281
rect -453 1281 -321 1297
rect -453 1264 -437 1281
rect -595 1247 -545 1264
rect -745 1200 -545 1247
rect -487 1247 -437 1264
rect -337 1264 -321 1281
rect -195 1281 -63 1297
rect -195 1264 -179 1281
rect -337 1247 -287 1264
rect -487 1200 -287 1247
rect -229 1247 -179 1264
rect -79 1264 -63 1281
rect 63 1281 195 1297
rect 63 1264 79 1281
rect -79 1247 -29 1264
rect -229 1200 -29 1247
rect 29 1247 79 1264
rect 179 1264 195 1281
rect 321 1281 453 1297
rect 321 1264 337 1281
rect 179 1247 229 1264
rect 29 1200 229 1247
rect 287 1247 337 1264
rect 437 1264 453 1281
rect 579 1281 711 1297
rect 579 1264 595 1281
rect 437 1247 487 1264
rect 287 1200 487 1247
rect 545 1247 595 1264
rect 695 1264 711 1281
rect 837 1281 969 1297
rect 837 1264 853 1281
rect 695 1247 745 1264
rect 545 1200 745 1247
rect 803 1247 853 1264
rect 953 1264 969 1281
rect 1095 1281 1227 1297
rect 1095 1264 1111 1281
rect 953 1247 1003 1264
rect 803 1200 1003 1247
rect 1061 1247 1111 1264
rect 1211 1264 1227 1281
rect 1353 1281 1485 1297
rect 1353 1264 1369 1281
rect 1211 1247 1261 1264
rect 1061 1200 1261 1247
rect 1319 1247 1369 1264
rect 1469 1264 1485 1281
rect 1611 1281 1743 1297
rect 1611 1264 1627 1281
rect 1469 1247 1519 1264
rect 1319 1200 1519 1247
rect 1577 1247 1627 1264
rect 1727 1264 1743 1281
rect 1869 1281 2001 1297
rect 1869 1264 1885 1281
rect 1727 1247 1777 1264
rect 1577 1200 1777 1247
rect 1835 1247 1885 1264
rect 1985 1264 2001 1281
rect 2127 1281 2259 1297
rect 2127 1264 2143 1281
rect 1985 1247 2035 1264
rect 1835 1200 2035 1247
rect 2093 1247 2143 1264
rect 2243 1264 2259 1281
rect 2385 1281 2517 1297
rect 2385 1264 2401 1281
rect 2243 1247 2293 1264
rect 2093 1200 2293 1247
rect 2351 1247 2401 1264
rect 2501 1264 2517 1281
rect 2643 1281 2775 1297
rect 2643 1264 2659 1281
rect 2501 1247 2551 1264
rect 2351 1200 2551 1247
rect 2609 1247 2659 1264
rect 2759 1264 2775 1281
rect 2901 1281 3033 1297
rect 2901 1264 2917 1281
rect 2759 1247 2809 1264
rect 2609 1200 2809 1247
rect 2867 1247 2917 1264
rect 3017 1264 3033 1281
rect 3159 1281 3291 1297
rect 3159 1264 3175 1281
rect 3017 1247 3067 1264
rect 2867 1200 3067 1247
rect 3125 1247 3175 1264
rect 3275 1264 3291 1281
rect 3417 1281 3549 1297
rect 3417 1264 3433 1281
rect 3275 1247 3325 1264
rect 3125 1200 3325 1247
rect 3383 1247 3433 1264
rect 3533 1264 3549 1281
rect 3675 1281 3807 1297
rect 3675 1264 3691 1281
rect 3533 1247 3583 1264
rect 3383 1200 3583 1247
rect 3641 1247 3691 1264
rect 3791 1264 3807 1281
rect 3933 1281 4065 1297
rect 3933 1264 3949 1281
rect 3791 1247 3841 1264
rect 3641 1200 3841 1247
rect 3899 1247 3949 1264
rect 4049 1264 4065 1281
rect 4191 1281 4323 1297
rect 4191 1264 4207 1281
rect 4049 1247 4099 1264
rect 3899 1200 4099 1247
rect 4157 1247 4207 1264
rect 4307 1264 4323 1281
rect 4449 1281 4581 1297
rect 4449 1264 4465 1281
rect 4307 1247 4357 1264
rect 4157 1200 4357 1247
rect 4415 1247 4465 1264
rect 4565 1264 4581 1281
rect 4707 1281 4839 1297
rect 4707 1264 4723 1281
rect 4565 1247 4615 1264
rect 4415 1200 4615 1247
rect 4673 1247 4723 1264
rect 4823 1264 4839 1281
rect 4965 1281 5097 1297
rect 4965 1264 4981 1281
rect 4823 1247 4873 1264
rect 4673 1200 4873 1247
rect 4931 1247 4981 1264
rect 5081 1264 5097 1281
rect 5081 1247 5131 1264
rect 4931 1200 5131 1247
rect -5131 -1247 -4931 -1200
rect -5131 -1264 -5081 -1247
rect -5097 -1281 -5081 -1264
rect -4981 -1264 -4931 -1247
rect -4873 -1247 -4673 -1200
rect -4873 -1264 -4823 -1247
rect -4981 -1281 -4965 -1264
rect -5097 -1297 -4965 -1281
rect -4839 -1281 -4823 -1264
rect -4723 -1264 -4673 -1247
rect -4615 -1247 -4415 -1200
rect -4615 -1264 -4565 -1247
rect -4723 -1281 -4707 -1264
rect -4839 -1297 -4707 -1281
rect -4581 -1281 -4565 -1264
rect -4465 -1264 -4415 -1247
rect -4357 -1247 -4157 -1200
rect -4357 -1264 -4307 -1247
rect -4465 -1281 -4449 -1264
rect -4581 -1297 -4449 -1281
rect -4323 -1281 -4307 -1264
rect -4207 -1264 -4157 -1247
rect -4099 -1247 -3899 -1200
rect -4099 -1264 -4049 -1247
rect -4207 -1281 -4191 -1264
rect -4323 -1297 -4191 -1281
rect -4065 -1281 -4049 -1264
rect -3949 -1264 -3899 -1247
rect -3841 -1247 -3641 -1200
rect -3841 -1264 -3791 -1247
rect -3949 -1281 -3933 -1264
rect -4065 -1297 -3933 -1281
rect -3807 -1281 -3791 -1264
rect -3691 -1264 -3641 -1247
rect -3583 -1247 -3383 -1200
rect -3583 -1264 -3533 -1247
rect -3691 -1281 -3675 -1264
rect -3807 -1297 -3675 -1281
rect -3549 -1281 -3533 -1264
rect -3433 -1264 -3383 -1247
rect -3325 -1247 -3125 -1200
rect -3325 -1264 -3275 -1247
rect -3433 -1281 -3417 -1264
rect -3549 -1297 -3417 -1281
rect -3291 -1281 -3275 -1264
rect -3175 -1264 -3125 -1247
rect -3067 -1247 -2867 -1200
rect -3067 -1264 -3017 -1247
rect -3175 -1281 -3159 -1264
rect -3291 -1297 -3159 -1281
rect -3033 -1281 -3017 -1264
rect -2917 -1264 -2867 -1247
rect -2809 -1247 -2609 -1200
rect -2809 -1264 -2759 -1247
rect -2917 -1281 -2901 -1264
rect -3033 -1297 -2901 -1281
rect -2775 -1281 -2759 -1264
rect -2659 -1264 -2609 -1247
rect -2551 -1247 -2351 -1200
rect -2551 -1264 -2501 -1247
rect -2659 -1281 -2643 -1264
rect -2775 -1297 -2643 -1281
rect -2517 -1281 -2501 -1264
rect -2401 -1264 -2351 -1247
rect -2293 -1247 -2093 -1200
rect -2293 -1264 -2243 -1247
rect -2401 -1281 -2385 -1264
rect -2517 -1297 -2385 -1281
rect -2259 -1281 -2243 -1264
rect -2143 -1264 -2093 -1247
rect -2035 -1247 -1835 -1200
rect -2035 -1264 -1985 -1247
rect -2143 -1281 -2127 -1264
rect -2259 -1297 -2127 -1281
rect -2001 -1281 -1985 -1264
rect -1885 -1264 -1835 -1247
rect -1777 -1247 -1577 -1200
rect -1777 -1264 -1727 -1247
rect -1885 -1281 -1869 -1264
rect -2001 -1297 -1869 -1281
rect -1743 -1281 -1727 -1264
rect -1627 -1264 -1577 -1247
rect -1519 -1247 -1319 -1200
rect -1519 -1264 -1469 -1247
rect -1627 -1281 -1611 -1264
rect -1743 -1297 -1611 -1281
rect -1485 -1281 -1469 -1264
rect -1369 -1264 -1319 -1247
rect -1261 -1247 -1061 -1200
rect -1261 -1264 -1211 -1247
rect -1369 -1281 -1353 -1264
rect -1485 -1297 -1353 -1281
rect -1227 -1281 -1211 -1264
rect -1111 -1264 -1061 -1247
rect -1003 -1247 -803 -1200
rect -1003 -1264 -953 -1247
rect -1111 -1281 -1095 -1264
rect -1227 -1297 -1095 -1281
rect -969 -1281 -953 -1264
rect -853 -1264 -803 -1247
rect -745 -1247 -545 -1200
rect -745 -1264 -695 -1247
rect -853 -1281 -837 -1264
rect -969 -1297 -837 -1281
rect -711 -1281 -695 -1264
rect -595 -1264 -545 -1247
rect -487 -1247 -287 -1200
rect -487 -1264 -437 -1247
rect -595 -1281 -579 -1264
rect -711 -1297 -579 -1281
rect -453 -1281 -437 -1264
rect -337 -1264 -287 -1247
rect -229 -1247 -29 -1200
rect -229 -1264 -179 -1247
rect -337 -1281 -321 -1264
rect -453 -1297 -321 -1281
rect -195 -1281 -179 -1264
rect -79 -1264 -29 -1247
rect 29 -1247 229 -1200
rect 29 -1264 79 -1247
rect -79 -1281 -63 -1264
rect -195 -1297 -63 -1281
rect 63 -1281 79 -1264
rect 179 -1264 229 -1247
rect 287 -1247 487 -1200
rect 287 -1264 337 -1247
rect 179 -1281 195 -1264
rect 63 -1297 195 -1281
rect 321 -1281 337 -1264
rect 437 -1264 487 -1247
rect 545 -1247 745 -1200
rect 545 -1264 595 -1247
rect 437 -1281 453 -1264
rect 321 -1297 453 -1281
rect 579 -1281 595 -1264
rect 695 -1264 745 -1247
rect 803 -1247 1003 -1200
rect 803 -1264 853 -1247
rect 695 -1281 711 -1264
rect 579 -1297 711 -1281
rect 837 -1281 853 -1264
rect 953 -1264 1003 -1247
rect 1061 -1247 1261 -1200
rect 1061 -1264 1111 -1247
rect 953 -1281 969 -1264
rect 837 -1297 969 -1281
rect 1095 -1281 1111 -1264
rect 1211 -1264 1261 -1247
rect 1319 -1247 1519 -1200
rect 1319 -1264 1369 -1247
rect 1211 -1281 1227 -1264
rect 1095 -1297 1227 -1281
rect 1353 -1281 1369 -1264
rect 1469 -1264 1519 -1247
rect 1577 -1247 1777 -1200
rect 1577 -1264 1627 -1247
rect 1469 -1281 1485 -1264
rect 1353 -1297 1485 -1281
rect 1611 -1281 1627 -1264
rect 1727 -1264 1777 -1247
rect 1835 -1247 2035 -1200
rect 1835 -1264 1885 -1247
rect 1727 -1281 1743 -1264
rect 1611 -1297 1743 -1281
rect 1869 -1281 1885 -1264
rect 1985 -1264 2035 -1247
rect 2093 -1247 2293 -1200
rect 2093 -1264 2143 -1247
rect 1985 -1281 2001 -1264
rect 1869 -1297 2001 -1281
rect 2127 -1281 2143 -1264
rect 2243 -1264 2293 -1247
rect 2351 -1247 2551 -1200
rect 2351 -1264 2401 -1247
rect 2243 -1281 2259 -1264
rect 2127 -1297 2259 -1281
rect 2385 -1281 2401 -1264
rect 2501 -1264 2551 -1247
rect 2609 -1247 2809 -1200
rect 2609 -1264 2659 -1247
rect 2501 -1281 2517 -1264
rect 2385 -1297 2517 -1281
rect 2643 -1281 2659 -1264
rect 2759 -1264 2809 -1247
rect 2867 -1247 3067 -1200
rect 2867 -1264 2917 -1247
rect 2759 -1281 2775 -1264
rect 2643 -1297 2775 -1281
rect 2901 -1281 2917 -1264
rect 3017 -1264 3067 -1247
rect 3125 -1247 3325 -1200
rect 3125 -1264 3175 -1247
rect 3017 -1281 3033 -1264
rect 2901 -1297 3033 -1281
rect 3159 -1281 3175 -1264
rect 3275 -1264 3325 -1247
rect 3383 -1247 3583 -1200
rect 3383 -1264 3433 -1247
rect 3275 -1281 3291 -1264
rect 3159 -1297 3291 -1281
rect 3417 -1281 3433 -1264
rect 3533 -1264 3583 -1247
rect 3641 -1247 3841 -1200
rect 3641 -1264 3691 -1247
rect 3533 -1281 3549 -1264
rect 3417 -1297 3549 -1281
rect 3675 -1281 3691 -1264
rect 3791 -1264 3841 -1247
rect 3899 -1247 4099 -1200
rect 3899 -1264 3949 -1247
rect 3791 -1281 3807 -1264
rect 3675 -1297 3807 -1281
rect 3933 -1281 3949 -1264
rect 4049 -1264 4099 -1247
rect 4157 -1247 4357 -1200
rect 4157 -1264 4207 -1247
rect 4049 -1281 4065 -1264
rect 3933 -1297 4065 -1281
rect 4191 -1281 4207 -1264
rect 4307 -1264 4357 -1247
rect 4415 -1247 4615 -1200
rect 4415 -1264 4465 -1247
rect 4307 -1281 4323 -1264
rect 4191 -1297 4323 -1281
rect 4449 -1281 4465 -1264
rect 4565 -1264 4615 -1247
rect 4673 -1247 4873 -1200
rect 4673 -1264 4723 -1247
rect 4565 -1281 4581 -1264
rect 4449 -1297 4581 -1281
rect 4707 -1281 4723 -1264
rect 4823 -1264 4873 -1247
rect 4931 -1247 5131 -1200
rect 4931 -1264 4981 -1247
rect 4823 -1281 4839 -1264
rect 4707 -1297 4839 -1281
rect 4965 -1281 4981 -1264
rect 5081 -1264 5131 -1247
rect 5081 -1281 5097 -1264
rect 4965 -1297 5097 -1281
<< polycont >>
rect -5081 1247 -4981 1281
rect -4823 1247 -4723 1281
rect -4565 1247 -4465 1281
rect -4307 1247 -4207 1281
rect -4049 1247 -3949 1281
rect -3791 1247 -3691 1281
rect -3533 1247 -3433 1281
rect -3275 1247 -3175 1281
rect -3017 1247 -2917 1281
rect -2759 1247 -2659 1281
rect -2501 1247 -2401 1281
rect -2243 1247 -2143 1281
rect -1985 1247 -1885 1281
rect -1727 1247 -1627 1281
rect -1469 1247 -1369 1281
rect -1211 1247 -1111 1281
rect -953 1247 -853 1281
rect -695 1247 -595 1281
rect -437 1247 -337 1281
rect -179 1247 -79 1281
rect 79 1247 179 1281
rect 337 1247 437 1281
rect 595 1247 695 1281
rect 853 1247 953 1281
rect 1111 1247 1211 1281
rect 1369 1247 1469 1281
rect 1627 1247 1727 1281
rect 1885 1247 1985 1281
rect 2143 1247 2243 1281
rect 2401 1247 2501 1281
rect 2659 1247 2759 1281
rect 2917 1247 3017 1281
rect 3175 1247 3275 1281
rect 3433 1247 3533 1281
rect 3691 1247 3791 1281
rect 3949 1247 4049 1281
rect 4207 1247 4307 1281
rect 4465 1247 4565 1281
rect 4723 1247 4823 1281
rect 4981 1247 5081 1281
rect -5081 -1281 -4981 -1247
rect -4823 -1281 -4723 -1247
rect -4565 -1281 -4465 -1247
rect -4307 -1281 -4207 -1247
rect -4049 -1281 -3949 -1247
rect -3791 -1281 -3691 -1247
rect -3533 -1281 -3433 -1247
rect -3275 -1281 -3175 -1247
rect -3017 -1281 -2917 -1247
rect -2759 -1281 -2659 -1247
rect -2501 -1281 -2401 -1247
rect -2243 -1281 -2143 -1247
rect -1985 -1281 -1885 -1247
rect -1727 -1281 -1627 -1247
rect -1469 -1281 -1369 -1247
rect -1211 -1281 -1111 -1247
rect -953 -1281 -853 -1247
rect -695 -1281 -595 -1247
rect -437 -1281 -337 -1247
rect -179 -1281 -79 -1247
rect 79 -1281 179 -1247
rect 337 -1281 437 -1247
rect 595 -1281 695 -1247
rect 853 -1281 953 -1247
rect 1111 -1281 1211 -1247
rect 1369 -1281 1469 -1247
rect 1627 -1281 1727 -1247
rect 1885 -1281 1985 -1247
rect 2143 -1281 2243 -1247
rect 2401 -1281 2501 -1247
rect 2659 -1281 2759 -1247
rect 2917 -1281 3017 -1247
rect 3175 -1281 3275 -1247
rect 3433 -1281 3533 -1247
rect 3691 -1281 3791 -1247
rect 3949 -1281 4049 -1247
rect 4207 -1281 4307 -1247
rect 4465 -1281 4565 -1247
rect 4723 -1281 4823 -1247
rect 4981 -1281 5081 -1247
<< locali >>
rect -5311 1385 -5215 1419
rect 5215 1385 5311 1419
rect -5311 1323 -5277 1385
rect 5277 1323 5311 1385
rect -5097 1247 -5081 1281
rect -4981 1247 -4965 1281
rect -4839 1247 -4823 1281
rect -4723 1247 -4707 1281
rect -4581 1247 -4565 1281
rect -4465 1247 -4449 1281
rect -4323 1247 -4307 1281
rect -4207 1247 -4191 1281
rect -4065 1247 -4049 1281
rect -3949 1247 -3933 1281
rect -3807 1247 -3791 1281
rect -3691 1247 -3675 1281
rect -3549 1247 -3533 1281
rect -3433 1247 -3417 1281
rect -3291 1247 -3275 1281
rect -3175 1247 -3159 1281
rect -3033 1247 -3017 1281
rect -2917 1247 -2901 1281
rect -2775 1247 -2759 1281
rect -2659 1247 -2643 1281
rect -2517 1247 -2501 1281
rect -2401 1247 -2385 1281
rect -2259 1247 -2243 1281
rect -2143 1247 -2127 1281
rect -2001 1247 -1985 1281
rect -1885 1247 -1869 1281
rect -1743 1247 -1727 1281
rect -1627 1247 -1611 1281
rect -1485 1247 -1469 1281
rect -1369 1247 -1353 1281
rect -1227 1247 -1211 1281
rect -1111 1247 -1095 1281
rect -969 1247 -953 1281
rect -853 1247 -837 1281
rect -711 1247 -695 1281
rect -595 1247 -579 1281
rect -453 1247 -437 1281
rect -337 1247 -321 1281
rect -195 1247 -179 1281
rect -79 1247 -63 1281
rect 63 1247 79 1281
rect 179 1247 195 1281
rect 321 1247 337 1281
rect 437 1247 453 1281
rect 579 1247 595 1281
rect 695 1247 711 1281
rect 837 1247 853 1281
rect 953 1247 969 1281
rect 1095 1247 1111 1281
rect 1211 1247 1227 1281
rect 1353 1247 1369 1281
rect 1469 1247 1485 1281
rect 1611 1247 1627 1281
rect 1727 1247 1743 1281
rect 1869 1247 1885 1281
rect 1985 1247 2001 1281
rect 2127 1247 2143 1281
rect 2243 1247 2259 1281
rect 2385 1247 2401 1281
rect 2501 1247 2517 1281
rect 2643 1247 2659 1281
rect 2759 1247 2775 1281
rect 2901 1247 2917 1281
rect 3017 1247 3033 1281
rect 3159 1247 3175 1281
rect 3275 1247 3291 1281
rect 3417 1247 3433 1281
rect 3533 1247 3549 1281
rect 3675 1247 3691 1281
rect 3791 1247 3807 1281
rect 3933 1247 3949 1281
rect 4049 1247 4065 1281
rect 4191 1247 4207 1281
rect 4307 1247 4323 1281
rect 4449 1247 4465 1281
rect 4565 1247 4581 1281
rect 4707 1247 4723 1281
rect 4823 1247 4839 1281
rect 4965 1247 4981 1281
rect 5081 1247 5097 1281
rect -5177 1188 -5143 1204
rect -5177 -1204 -5143 -1188
rect -4919 1188 -4885 1204
rect -4919 -1204 -4885 -1188
rect -4661 1188 -4627 1204
rect -4661 -1204 -4627 -1188
rect -4403 1188 -4369 1204
rect -4403 -1204 -4369 -1188
rect -4145 1188 -4111 1204
rect -4145 -1204 -4111 -1188
rect -3887 1188 -3853 1204
rect -3887 -1204 -3853 -1188
rect -3629 1188 -3595 1204
rect -3629 -1204 -3595 -1188
rect -3371 1188 -3337 1204
rect -3371 -1204 -3337 -1188
rect -3113 1188 -3079 1204
rect -3113 -1204 -3079 -1188
rect -2855 1188 -2821 1204
rect -2855 -1204 -2821 -1188
rect -2597 1188 -2563 1204
rect -2597 -1204 -2563 -1188
rect -2339 1188 -2305 1204
rect -2339 -1204 -2305 -1188
rect -2081 1188 -2047 1204
rect -2081 -1204 -2047 -1188
rect -1823 1188 -1789 1204
rect -1823 -1204 -1789 -1188
rect -1565 1188 -1531 1204
rect -1565 -1204 -1531 -1188
rect -1307 1188 -1273 1204
rect -1307 -1204 -1273 -1188
rect -1049 1188 -1015 1204
rect -1049 -1204 -1015 -1188
rect -791 1188 -757 1204
rect -791 -1204 -757 -1188
rect -533 1188 -499 1204
rect -533 -1204 -499 -1188
rect -275 1188 -241 1204
rect -275 -1204 -241 -1188
rect -17 1188 17 1204
rect -17 -1204 17 -1188
rect 241 1188 275 1204
rect 241 -1204 275 -1188
rect 499 1188 533 1204
rect 499 -1204 533 -1188
rect 757 1188 791 1204
rect 757 -1204 791 -1188
rect 1015 1188 1049 1204
rect 1015 -1204 1049 -1188
rect 1273 1188 1307 1204
rect 1273 -1204 1307 -1188
rect 1531 1188 1565 1204
rect 1531 -1204 1565 -1188
rect 1789 1188 1823 1204
rect 1789 -1204 1823 -1188
rect 2047 1188 2081 1204
rect 2047 -1204 2081 -1188
rect 2305 1188 2339 1204
rect 2305 -1204 2339 -1188
rect 2563 1188 2597 1204
rect 2563 -1204 2597 -1188
rect 2821 1188 2855 1204
rect 2821 -1204 2855 -1188
rect 3079 1188 3113 1204
rect 3079 -1204 3113 -1188
rect 3337 1188 3371 1204
rect 3337 -1204 3371 -1188
rect 3595 1188 3629 1204
rect 3595 -1204 3629 -1188
rect 3853 1188 3887 1204
rect 3853 -1204 3887 -1188
rect 4111 1188 4145 1204
rect 4111 -1204 4145 -1188
rect 4369 1188 4403 1204
rect 4369 -1204 4403 -1188
rect 4627 1188 4661 1204
rect 4627 -1204 4661 -1188
rect 4885 1188 4919 1204
rect 4885 -1204 4919 -1188
rect 5143 1188 5177 1204
rect 5143 -1204 5177 -1188
rect -5097 -1281 -5081 -1247
rect -4981 -1281 -4965 -1247
rect -4839 -1281 -4823 -1247
rect -4723 -1281 -4707 -1247
rect -4581 -1281 -4565 -1247
rect -4465 -1281 -4449 -1247
rect -4323 -1281 -4307 -1247
rect -4207 -1281 -4191 -1247
rect -4065 -1281 -4049 -1247
rect -3949 -1281 -3933 -1247
rect -3807 -1281 -3791 -1247
rect -3691 -1281 -3675 -1247
rect -3549 -1281 -3533 -1247
rect -3433 -1281 -3417 -1247
rect -3291 -1281 -3275 -1247
rect -3175 -1281 -3159 -1247
rect -3033 -1281 -3017 -1247
rect -2917 -1281 -2901 -1247
rect -2775 -1281 -2759 -1247
rect -2659 -1281 -2643 -1247
rect -2517 -1281 -2501 -1247
rect -2401 -1281 -2385 -1247
rect -2259 -1281 -2243 -1247
rect -2143 -1281 -2127 -1247
rect -2001 -1281 -1985 -1247
rect -1885 -1281 -1869 -1247
rect -1743 -1281 -1727 -1247
rect -1627 -1281 -1611 -1247
rect -1485 -1281 -1469 -1247
rect -1369 -1281 -1353 -1247
rect -1227 -1281 -1211 -1247
rect -1111 -1281 -1095 -1247
rect -969 -1281 -953 -1247
rect -853 -1281 -837 -1247
rect -711 -1281 -695 -1247
rect -595 -1281 -579 -1247
rect -453 -1281 -437 -1247
rect -337 -1281 -321 -1247
rect -195 -1281 -179 -1247
rect -79 -1281 -63 -1247
rect 63 -1281 79 -1247
rect 179 -1281 195 -1247
rect 321 -1281 337 -1247
rect 437 -1281 453 -1247
rect 579 -1281 595 -1247
rect 695 -1281 711 -1247
rect 837 -1281 853 -1247
rect 953 -1281 969 -1247
rect 1095 -1281 1111 -1247
rect 1211 -1281 1227 -1247
rect 1353 -1281 1369 -1247
rect 1469 -1281 1485 -1247
rect 1611 -1281 1627 -1247
rect 1727 -1281 1743 -1247
rect 1869 -1281 1885 -1247
rect 1985 -1281 2001 -1247
rect 2127 -1281 2143 -1247
rect 2243 -1281 2259 -1247
rect 2385 -1281 2401 -1247
rect 2501 -1281 2517 -1247
rect 2643 -1281 2659 -1247
rect 2759 -1281 2775 -1247
rect 2901 -1281 2917 -1247
rect 3017 -1281 3033 -1247
rect 3159 -1281 3175 -1247
rect 3275 -1281 3291 -1247
rect 3417 -1281 3433 -1247
rect 3533 -1281 3549 -1247
rect 3675 -1281 3691 -1247
rect 3791 -1281 3807 -1247
rect 3933 -1281 3949 -1247
rect 4049 -1281 4065 -1247
rect 4191 -1281 4207 -1247
rect 4307 -1281 4323 -1247
rect 4449 -1281 4465 -1247
rect 4565 -1281 4581 -1247
rect 4707 -1281 4723 -1247
rect 4823 -1281 4839 -1247
rect 4965 -1281 4981 -1247
rect 5081 -1281 5097 -1247
rect -5311 -1385 -5277 -1323
rect 5277 -1385 5311 -1323
rect -5311 -1419 -5215 -1385
rect 5215 -1419 5311 -1385
<< viali >>
rect -5081 1247 -4981 1281
rect -4823 1247 -4723 1281
rect -4565 1247 -4465 1281
rect -4307 1247 -4207 1281
rect -4049 1247 -3949 1281
rect -3791 1247 -3691 1281
rect -3533 1247 -3433 1281
rect -3275 1247 -3175 1281
rect -3017 1247 -2917 1281
rect -2759 1247 -2659 1281
rect -2501 1247 -2401 1281
rect -2243 1247 -2143 1281
rect -1985 1247 -1885 1281
rect -1727 1247 -1627 1281
rect -1469 1247 -1369 1281
rect -1211 1247 -1111 1281
rect -953 1247 -853 1281
rect -695 1247 -595 1281
rect -437 1247 -337 1281
rect -179 1247 -79 1281
rect 79 1247 179 1281
rect 337 1247 437 1281
rect 595 1247 695 1281
rect 853 1247 953 1281
rect 1111 1247 1211 1281
rect 1369 1247 1469 1281
rect 1627 1247 1727 1281
rect 1885 1247 1985 1281
rect 2143 1247 2243 1281
rect 2401 1247 2501 1281
rect 2659 1247 2759 1281
rect 2917 1247 3017 1281
rect 3175 1247 3275 1281
rect 3433 1247 3533 1281
rect 3691 1247 3791 1281
rect 3949 1247 4049 1281
rect 4207 1247 4307 1281
rect 4465 1247 4565 1281
rect 4723 1247 4823 1281
rect 4981 1247 5081 1281
rect -5177 -1188 -5143 1188
rect -4919 -1188 -4885 1188
rect -4661 -1188 -4627 1188
rect -4403 -1188 -4369 1188
rect -4145 -1188 -4111 1188
rect -3887 -1188 -3853 1188
rect -3629 -1188 -3595 1188
rect -3371 -1188 -3337 1188
rect -3113 -1188 -3079 1188
rect -2855 -1188 -2821 1188
rect -2597 -1188 -2563 1188
rect -2339 -1188 -2305 1188
rect -2081 -1188 -2047 1188
rect -1823 -1188 -1789 1188
rect -1565 -1188 -1531 1188
rect -1307 -1188 -1273 1188
rect -1049 -1188 -1015 1188
rect -791 -1188 -757 1188
rect -533 -1188 -499 1188
rect -275 -1188 -241 1188
rect -17 -1188 17 1188
rect 241 -1188 275 1188
rect 499 -1188 533 1188
rect 757 -1188 791 1188
rect 1015 -1188 1049 1188
rect 1273 -1188 1307 1188
rect 1531 -1188 1565 1188
rect 1789 -1188 1823 1188
rect 2047 -1188 2081 1188
rect 2305 -1188 2339 1188
rect 2563 -1188 2597 1188
rect 2821 -1188 2855 1188
rect 3079 -1188 3113 1188
rect 3337 -1188 3371 1188
rect 3595 -1188 3629 1188
rect 3853 -1188 3887 1188
rect 4111 -1188 4145 1188
rect 4369 -1188 4403 1188
rect 4627 -1188 4661 1188
rect 4885 -1188 4919 1188
rect 5143 -1188 5177 1188
rect -5081 -1281 -4981 -1247
rect -4823 -1281 -4723 -1247
rect -4565 -1281 -4465 -1247
rect -4307 -1281 -4207 -1247
rect -4049 -1281 -3949 -1247
rect -3791 -1281 -3691 -1247
rect -3533 -1281 -3433 -1247
rect -3275 -1281 -3175 -1247
rect -3017 -1281 -2917 -1247
rect -2759 -1281 -2659 -1247
rect -2501 -1281 -2401 -1247
rect -2243 -1281 -2143 -1247
rect -1985 -1281 -1885 -1247
rect -1727 -1281 -1627 -1247
rect -1469 -1281 -1369 -1247
rect -1211 -1281 -1111 -1247
rect -953 -1281 -853 -1247
rect -695 -1281 -595 -1247
rect -437 -1281 -337 -1247
rect -179 -1281 -79 -1247
rect 79 -1281 179 -1247
rect 337 -1281 437 -1247
rect 595 -1281 695 -1247
rect 853 -1281 953 -1247
rect 1111 -1281 1211 -1247
rect 1369 -1281 1469 -1247
rect 1627 -1281 1727 -1247
rect 1885 -1281 1985 -1247
rect 2143 -1281 2243 -1247
rect 2401 -1281 2501 -1247
rect 2659 -1281 2759 -1247
rect 2917 -1281 3017 -1247
rect 3175 -1281 3275 -1247
rect 3433 -1281 3533 -1247
rect 3691 -1281 3791 -1247
rect 3949 -1281 4049 -1247
rect 4207 -1281 4307 -1247
rect 4465 -1281 4565 -1247
rect 4723 -1281 4823 -1247
rect 4981 -1281 5081 -1247
<< metal1 >>
rect -5093 1281 -4969 1287
rect -5093 1247 -5081 1281
rect -4981 1247 -4969 1281
rect -5093 1241 -4969 1247
rect -4835 1281 -4711 1287
rect -4835 1247 -4823 1281
rect -4723 1247 -4711 1281
rect -4835 1241 -4711 1247
rect -4577 1281 -4453 1287
rect -4577 1247 -4565 1281
rect -4465 1247 -4453 1281
rect -4577 1241 -4453 1247
rect -4319 1281 -4195 1287
rect -4319 1247 -4307 1281
rect -4207 1247 -4195 1281
rect -4319 1241 -4195 1247
rect -4061 1281 -3937 1287
rect -4061 1247 -4049 1281
rect -3949 1247 -3937 1281
rect -4061 1241 -3937 1247
rect -3803 1281 -3679 1287
rect -3803 1247 -3791 1281
rect -3691 1247 -3679 1281
rect -3803 1241 -3679 1247
rect -3545 1281 -3421 1287
rect -3545 1247 -3533 1281
rect -3433 1247 -3421 1281
rect -3545 1241 -3421 1247
rect -3287 1281 -3163 1287
rect -3287 1247 -3275 1281
rect -3175 1247 -3163 1281
rect -3287 1241 -3163 1247
rect -3029 1281 -2905 1287
rect -3029 1247 -3017 1281
rect -2917 1247 -2905 1281
rect -3029 1241 -2905 1247
rect -2771 1281 -2647 1287
rect -2771 1247 -2759 1281
rect -2659 1247 -2647 1281
rect -2771 1241 -2647 1247
rect -2513 1281 -2389 1287
rect -2513 1247 -2501 1281
rect -2401 1247 -2389 1281
rect -2513 1241 -2389 1247
rect -2255 1281 -2131 1287
rect -2255 1247 -2243 1281
rect -2143 1247 -2131 1281
rect -2255 1241 -2131 1247
rect -1997 1281 -1873 1287
rect -1997 1247 -1985 1281
rect -1885 1247 -1873 1281
rect -1997 1241 -1873 1247
rect -1739 1281 -1615 1287
rect -1739 1247 -1727 1281
rect -1627 1247 -1615 1281
rect -1739 1241 -1615 1247
rect -1481 1281 -1357 1287
rect -1481 1247 -1469 1281
rect -1369 1247 -1357 1281
rect -1481 1241 -1357 1247
rect -1223 1281 -1099 1287
rect -1223 1247 -1211 1281
rect -1111 1247 -1099 1281
rect -1223 1241 -1099 1247
rect -965 1281 -841 1287
rect -965 1247 -953 1281
rect -853 1247 -841 1281
rect -965 1241 -841 1247
rect -707 1281 -583 1287
rect -707 1247 -695 1281
rect -595 1247 -583 1281
rect -707 1241 -583 1247
rect -449 1281 -325 1287
rect -449 1247 -437 1281
rect -337 1247 -325 1281
rect -449 1241 -325 1247
rect -191 1281 -67 1287
rect -191 1247 -179 1281
rect -79 1247 -67 1281
rect -191 1241 -67 1247
rect 67 1281 191 1287
rect 67 1247 79 1281
rect 179 1247 191 1281
rect 67 1241 191 1247
rect 325 1281 449 1287
rect 325 1247 337 1281
rect 437 1247 449 1281
rect 325 1241 449 1247
rect 583 1281 707 1287
rect 583 1247 595 1281
rect 695 1247 707 1281
rect 583 1241 707 1247
rect 841 1281 965 1287
rect 841 1247 853 1281
rect 953 1247 965 1281
rect 841 1241 965 1247
rect 1099 1281 1223 1287
rect 1099 1247 1111 1281
rect 1211 1247 1223 1281
rect 1099 1241 1223 1247
rect 1357 1281 1481 1287
rect 1357 1247 1369 1281
rect 1469 1247 1481 1281
rect 1357 1241 1481 1247
rect 1615 1281 1739 1287
rect 1615 1247 1627 1281
rect 1727 1247 1739 1281
rect 1615 1241 1739 1247
rect 1873 1281 1997 1287
rect 1873 1247 1885 1281
rect 1985 1247 1997 1281
rect 1873 1241 1997 1247
rect 2131 1281 2255 1287
rect 2131 1247 2143 1281
rect 2243 1247 2255 1281
rect 2131 1241 2255 1247
rect 2389 1281 2513 1287
rect 2389 1247 2401 1281
rect 2501 1247 2513 1281
rect 2389 1241 2513 1247
rect 2647 1281 2771 1287
rect 2647 1247 2659 1281
rect 2759 1247 2771 1281
rect 2647 1241 2771 1247
rect 2905 1281 3029 1287
rect 2905 1247 2917 1281
rect 3017 1247 3029 1281
rect 2905 1241 3029 1247
rect 3163 1281 3287 1287
rect 3163 1247 3175 1281
rect 3275 1247 3287 1281
rect 3163 1241 3287 1247
rect 3421 1281 3545 1287
rect 3421 1247 3433 1281
rect 3533 1247 3545 1281
rect 3421 1241 3545 1247
rect 3679 1281 3803 1287
rect 3679 1247 3691 1281
rect 3791 1247 3803 1281
rect 3679 1241 3803 1247
rect 3937 1281 4061 1287
rect 3937 1247 3949 1281
rect 4049 1247 4061 1281
rect 3937 1241 4061 1247
rect 4195 1281 4319 1287
rect 4195 1247 4207 1281
rect 4307 1247 4319 1281
rect 4195 1241 4319 1247
rect 4453 1281 4577 1287
rect 4453 1247 4465 1281
rect 4565 1247 4577 1281
rect 4453 1241 4577 1247
rect 4711 1281 4835 1287
rect 4711 1247 4723 1281
rect 4823 1247 4835 1281
rect 4711 1241 4835 1247
rect 4969 1281 5093 1287
rect 4969 1247 4981 1281
rect 5081 1247 5093 1281
rect 4969 1241 5093 1247
rect -5183 1188 -5137 1200
rect -5183 -1188 -5177 1188
rect -5143 -1188 -5137 1188
rect -5183 -1200 -5137 -1188
rect -4925 1188 -4879 1200
rect -4925 -1188 -4919 1188
rect -4885 -1188 -4879 1188
rect -4925 -1200 -4879 -1188
rect -4667 1188 -4621 1200
rect -4667 -1188 -4661 1188
rect -4627 -1188 -4621 1188
rect -4667 -1200 -4621 -1188
rect -4409 1188 -4363 1200
rect -4409 -1188 -4403 1188
rect -4369 -1188 -4363 1188
rect -4409 -1200 -4363 -1188
rect -4151 1188 -4105 1200
rect -4151 -1188 -4145 1188
rect -4111 -1188 -4105 1188
rect -4151 -1200 -4105 -1188
rect -3893 1188 -3847 1200
rect -3893 -1188 -3887 1188
rect -3853 -1188 -3847 1188
rect -3893 -1200 -3847 -1188
rect -3635 1188 -3589 1200
rect -3635 -1188 -3629 1188
rect -3595 -1188 -3589 1188
rect -3635 -1200 -3589 -1188
rect -3377 1188 -3331 1200
rect -3377 -1188 -3371 1188
rect -3337 -1188 -3331 1188
rect -3377 -1200 -3331 -1188
rect -3119 1188 -3073 1200
rect -3119 -1188 -3113 1188
rect -3079 -1188 -3073 1188
rect -3119 -1200 -3073 -1188
rect -2861 1188 -2815 1200
rect -2861 -1188 -2855 1188
rect -2821 -1188 -2815 1188
rect -2861 -1200 -2815 -1188
rect -2603 1188 -2557 1200
rect -2603 -1188 -2597 1188
rect -2563 -1188 -2557 1188
rect -2603 -1200 -2557 -1188
rect -2345 1188 -2299 1200
rect -2345 -1188 -2339 1188
rect -2305 -1188 -2299 1188
rect -2345 -1200 -2299 -1188
rect -2087 1188 -2041 1200
rect -2087 -1188 -2081 1188
rect -2047 -1188 -2041 1188
rect -2087 -1200 -2041 -1188
rect -1829 1188 -1783 1200
rect -1829 -1188 -1823 1188
rect -1789 -1188 -1783 1188
rect -1829 -1200 -1783 -1188
rect -1571 1188 -1525 1200
rect -1571 -1188 -1565 1188
rect -1531 -1188 -1525 1188
rect -1571 -1200 -1525 -1188
rect -1313 1188 -1267 1200
rect -1313 -1188 -1307 1188
rect -1273 -1188 -1267 1188
rect -1313 -1200 -1267 -1188
rect -1055 1188 -1009 1200
rect -1055 -1188 -1049 1188
rect -1015 -1188 -1009 1188
rect -1055 -1200 -1009 -1188
rect -797 1188 -751 1200
rect -797 -1188 -791 1188
rect -757 -1188 -751 1188
rect -797 -1200 -751 -1188
rect -539 1188 -493 1200
rect -539 -1188 -533 1188
rect -499 -1188 -493 1188
rect -539 -1200 -493 -1188
rect -281 1188 -235 1200
rect -281 -1188 -275 1188
rect -241 -1188 -235 1188
rect -281 -1200 -235 -1188
rect -23 1188 23 1200
rect -23 -1188 -17 1188
rect 17 -1188 23 1188
rect -23 -1200 23 -1188
rect 235 1188 281 1200
rect 235 -1188 241 1188
rect 275 -1188 281 1188
rect 235 -1200 281 -1188
rect 493 1188 539 1200
rect 493 -1188 499 1188
rect 533 -1188 539 1188
rect 493 -1200 539 -1188
rect 751 1188 797 1200
rect 751 -1188 757 1188
rect 791 -1188 797 1188
rect 751 -1200 797 -1188
rect 1009 1188 1055 1200
rect 1009 -1188 1015 1188
rect 1049 -1188 1055 1188
rect 1009 -1200 1055 -1188
rect 1267 1188 1313 1200
rect 1267 -1188 1273 1188
rect 1307 -1188 1313 1188
rect 1267 -1200 1313 -1188
rect 1525 1188 1571 1200
rect 1525 -1188 1531 1188
rect 1565 -1188 1571 1188
rect 1525 -1200 1571 -1188
rect 1783 1188 1829 1200
rect 1783 -1188 1789 1188
rect 1823 -1188 1829 1188
rect 1783 -1200 1829 -1188
rect 2041 1188 2087 1200
rect 2041 -1188 2047 1188
rect 2081 -1188 2087 1188
rect 2041 -1200 2087 -1188
rect 2299 1188 2345 1200
rect 2299 -1188 2305 1188
rect 2339 -1188 2345 1188
rect 2299 -1200 2345 -1188
rect 2557 1188 2603 1200
rect 2557 -1188 2563 1188
rect 2597 -1188 2603 1188
rect 2557 -1200 2603 -1188
rect 2815 1188 2861 1200
rect 2815 -1188 2821 1188
rect 2855 -1188 2861 1188
rect 2815 -1200 2861 -1188
rect 3073 1188 3119 1200
rect 3073 -1188 3079 1188
rect 3113 -1188 3119 1188
rect 3073 -1200 3119 -1188
rect 3331 1188 3377 1200
rect 3331 -1188 3337 1188
rect 3371 -1188 3377 1188
rect 3331 -1200 3377 -1188
rect 3589 1188 3635 1200
rect 3589 -1188 3595 1188
rect 3629 -1188 3635 1188
rect 3589 -1200 3635 -1188
rect 3847 1188 3893 1200
rect 3847 -1188 3853 1188
rect 3887 -1188 3893 1188
rect 3847 -1200 3893 -1188
rect 4105 1188 4151 1200
rect 4105 -1188 4111 1188
rect 4145 -1188 4151 1188
rect 4105 -1200 4151 -1188
rect 4363 1188 4409 1200
rect 4363 -1188 4369 1188
rect 4403 -1188 4409 1188
rect 4363 -1200 4409 -1188
rect 4621 1188 4667 1200
rect 4621 -1188 4627 1188
rect 4661 -1188 4667 1188
rect 4621 -1200 4667 -1188
rect 4879 1188 4925 1200
rect 4879 -1188 4885 1188
rect 4919 -1188 4925 1188
rect 4879 -1200 4925 -1188
rect 5137 1188 5183 1200
rect 5137 -1188 5143 1188
rect 5177 -1188 5183 1188
rect 5137 -1200 5183 -1188
rect -5093 -1247 -4969 -1241
rect -5093 -1281 -5081 -1247
rect -4981 -1281 -4969 -1247
rect -5093 -1287 -4969 -1281
rect -4835 -1247 -4711 -1241
rect -4835 -1281 -4823 -1247
rect -4723 -1281 -4711 -1247
rect -4835 -1287 -4711 -1281
rect -4577 -1247 -4453 -1241
rect -4577 -1281 -4565 -1247
rect -4465 -1281 -4453 -1247
rect -4577 -1287 -4453 -1281
rect -4319 -1247 -4195 -1241
rect -4319 -1281 -4307 -1247
rect -4207 -1281 -4195 -1247
rect -4319 -1287 -4195 -1281
rect -4061 -1247 -3937 -1241
rect -4061 -1281 -4049 -1247
rect -3949 -1281 -3937 -1247
rect -4061 -1287 -3937 -1281
rect -3803 -1247 -3679 -1241
rect -3803 -1281 -3791 -1247
rect -3691 -1281 -3679 -1247
rect -3803 -1287 -3679 -1281
rect -3545 -1247 -3421 -1241
rect -3545 -1281 -3533 -1247
rect -3433 -1281 -3421 -1247
rect -3545 -1287 -3421 -1281
rect -3287 -1247 -3163 -1241
rect -3287 -1281 -3275 -1247
rect -3175 -1281 -3163 -1247
rect -3287 -1287 -3163 -1281
rect -3029 -1247 -2905 -1241
rect -3029 -1281 -3017 -1247
rect -2917 -1281 -2905 -1247
rect -3029 -1287 -2905 -1281
rect -2771 -1247 -2647 -1241
rect -2771 -1281 -2759 -1247
rect -2659 -1281 -2647 -1247
rect -2771 -1287 -2647 -1281
rect -2513 -1247 -2389 -1241
rect -2513 -1281 -2501 -1247
rect -2401 -1281 -2389 -1247
rect -2513 -1287 -2389 -1281
rect -2255 -1247 -2131 -1241
rect -2255 -1281 -2243 -1247
rect -2143 -1281 -2131 -1247
rect -2255 -1287 -2131 -1281
rect -1997 -1247 -1873 -1241
rect -1997 -1281 -1985 -1247
rect -1885 -1281 -1873 -1247
rect -1997 -1287 -1873 -1281
rect -1739 -1247 -1615 -1241
rect -1739 -1281 -1727 -1247
rect -1627 -1281 -1615 -1247
rect -1739 -1287 -1615 -1281
rect -1481 -1247 -1357 -1241
rect -1481 -1281 -1469 -1247
rect -1369 -1281 -1357 -1247
rect -1481 -1287 -1357 -1281
rect -1223 -1247 -1099 -1241
rect -1223 -1281 -1211 -1247
rect -1111 -1281 -1099 -1247
rect -1223 -1287 -1099 -1281
rect -965 -1247 -841 -1241
rect -965 -1281 -953 -1247
rect -853 -1281 -841 -1247
rect -965 -1287 -841 -1281
rect -707 -1247 -583 -1241
rect -707 -1281 -695 -1247
rect -595 -1281 -583 -1247
rect -707 -1287 -583 -1281
rect -449 -1247 -325 -1241
rect -449 -1281 -437 -1247
rect -337 -1281 -325 -1247
rect -449 -1287 -325 -1281
rect -191 -1247 -67 -1241
rect -191 -1281 -179 -1247
rect -79 -1281 -67 -1247
rect -191 -1287 -67 -1281
rect 67 -1247 191 -1241
rect 67 -1281 79 -1247
rect 179 -1281 191 -1247
rect 67 -1287 191 -1281
rect 325 -1247 449 -1241
rect 325 -1281 337 -1247
rect 437 -1281 449 -1247
rect 325 -1287 449 -1281
rect 583 -1247 707 -1241
rect 583 -1281 595 -1247
rect 695 -1281 707 -1247
rect 583 -1287 707 -1281
rect 841 -1247 965 -1241
rect 841 -1281 853 -1247
rect 953 -1281 965 -1247
rect 841 -1287 965 -1281
rect 1099 -1247 1223 -1241
rect 1099 -1281 1111 -1247
rect 1211 -1281 1223 -1247
rect 1099 -1287 1223 -1281
rect 1357 -1247 1481 -1241
rect 1357 -1281 1369 -1247
rect 1469 -1281 1481 -1247
rect 1357 -1287 1481 -1281
rect 1615 -1247 1739 -1241
rect 1615 -1281 1627 -1247
rect 1727 -1281 1739 -1247
rect 1615 -1287 1739 -1281
rect 1873 -1247 1997 -1241
rect 1873 -1281 1885 -1247
rect 1985 -1281 1997 -1247
rect 1873 -1287 1997 -1281
rect 2131 -1247 2255 -1241
rect 2131 -1281 2143 -1247
rect 2243 -1281 2255 -1247
rect 2131 -1287 2255 -1281
rect 2389 -1247 2513 -1241
rect 2389 -1281 2401 -1247
rect 2501 -1281 2513 -1247
rect 2389 -1287 2513 -1281
rect 2647 -1247 2771 -1241
rect 2647 -1281 2659 -1247
rect 2759 -1281 2771 -1247
rect 2647 -1287 2771 -1281
rect 2905 -1247 3029 -1241
rect 2905 -1281 2917 -1247
rect 3017 -1281 3029 -1247
rect 2905 -1287 3029 -1281
rect 3163 -1247 3287 -1241
rect 3163 -1281 3175 -1247
rect 3275 -1281 3287 -1247
rect 3163 -1287 3287 -1281
rect 3421 -1247 3545 -1241
rect 3421 -1281 3433 -1247
rect 3533 -1281 3545 -1247
rect 3421 -1287 3545 -1281
rect 3679 -1247 3803 -1241
rect 3679 -1281 3691 -1247
rect 3791 -1281 3803 -1247
rect 3679 -1287 3803 -1281
rect 3937 -1247 4061 -1241
rect 3937 -1281 3949 -1247
rect 4049 -1281 4061 -1247
rect 3937 -1287 4061 -1281
rect 4195 -1247 4319 -1241
rect 4195 -1281 4207 -1247
rect 4307 -1281 4319 -1247
rect 4195 -1287 4319 -1281
rect 4453 -1247 4577 -1241
rect 4453 -1281 4465 -1247
rect 4565 -1281 4577 -1247
rect 4453 -1287 4577 -1281
rect 4711 -1247 4835 -1241
rect 4711 -1281 4723 -1247
rect 4823 -1281 4835 -1247
rect 4711 -1287 4835 -1281
rect 4969 -1247 5093 -1241
rect 4969 -1281 4981 -1247
rect 5081 -1281 5093 -1247
rect 4969 -1287 5093 -1281
<< properties >>
string FIXED_BBOX -5294 -1402 5294 1402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 12 l 1 m 1 nf 40 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713232886
<< pwell >>
rect -2521 -2367 2521 2367
<< mvnmos >>
rect -2293 109 -2093 2109
rect -2035 109 -1835 2109
rect -1777 109 -1577 2109
rect -1519 109 -1319 2109
rect -1261 109 -1061 2109
rect -1003 109 -803 2109
rect -745 109 -545 2109
rect -487 109 -287 2109
rect -229 109 -29 2109
rect 29 109 229 2109
rect 287 109 487 2109
rect 545 109 745 2109
rect 803 109 1003 2109
rect 1061 109 1261 2109
rect 1319 109 1519 2109
rect 1577 109 1777 2109
rect 1835 109 2035 2109
rect 2093 109 2293 2109
rect -2293 -2109 -2093 -109
rect -2035 -2109 -1835 -109
rect -1777 -2109 -1577 -109
rect -1519 -2109 -1319 -109
rect -1261 -2109 -1061 -109
rect -1003 -2109 -803 -109
rect -745 -2109 -545 -109
rect -487 -2109 -287 -109
rect -229 -2109 -29 -109
rect 29 -2109 229 -109
rect 287 -2109 487 -109
rect 545 -2109 745 -109
rect 803 -2109 1003 -109
rect 1061 -2109 1261 -109
rect 1319 -2109 1519 -109
rect 1577 -2109 1777 -109
rect 1835 -2109 2035 -109
rect 2093 -2109 2293 -109
<< mvndiff >>
rect -2351 2097 -2293 2109
rect -2351 121 -2339 2097
rect -2305 121 -2293 2097
rect -2351 109 -2293 121
rect -2093 2097 -2035 2109
rect -2093 121 -2081 2097
rect -2047 121 -2035 2097
rect -2093 109 -2035 121
rect -1835 2097 -1777 2109
rect -1835 121 -1823 2097
rect -1789 121 -1777 2097
rect -1835 109 -1777 121
rect -1577 2097 -1519 2109
rect -1577 121 -1565 2097
rect -1531 121 -1519 2097
rect -1577 109 -1519 121
rect -1319 2097 -1261 2109
rect -1319 121 -1307 2097
rect -1273 121 -1261 2097
rect -1319 109 -1261 121
rect -1061 2097 -1003 2109
rect -1061 121 -1049 2097
rect -1015 121 -1003 2097
rect -1061 109 -1003 121
rect -803 2097 -745 2109
rect -803 121 -791 2097
rect -757 121 -745 2097
rect -803 109 -745 121
rect -545 2097 -487 2109
rect -545 121 -533 2097
rect -499 121 -487 2097
rect -545 109 -487 121
rect -287 2097 -229 2109
rect -287 121 -275 2097
rect -241 121 -229 2097
rect -287 109 -229 121
rect -29 2097 29 2109
rect -29 121 -17 2097
rect 17 121 29 2097
rect -29 109 29 121
rect 229 2097 287 2109
rect 229 121 241 2097
rect 275 121 287 2097
rect 229 109 287 121
rect 487 2097 545 2109
rect 487 121 499 2097
rect 533 121 545 2097
rect 487 109 545 121
rect 745 2097 803 2109
rect 745 121 757 2097
rect 791 121 803 2097
rect 745 109 803 121
rect 1003 2097 1061 2109
rect 1003 121 1015 2097
rect 1049 121 1061 2097
rect 1003 109 1061 121
rect 1261 2097 1319 2109
rect 1261 121 1273 2097
rect 1307 121 1319 2097
rect 1261 109 1319 121
rect 1519 2097 1577 2109
rect 1519 121 1531 2097
rect 1565 121 1577 2097
rect 1519 109 1577 121
rect 1777 2097 1835 2109
rect 1777 121 1789 2097
rect 1823 121 1835 2097
rect 1777 109 1835 121
rect 2035 2097 2093 2109
rect 2035 121 2047 2097
rect 2081 121 2093 2097
rect 2035 109 2093 121
rect 2293 2097 2351 2109
rect 2293 121 2305 2097
rect 2339 121 2351 2097
rect 2293 109 2351 121
rect -2351 -121 -2293 -109
rect -2351 -2097 -2339 -121
rect -2305 -2097 -2293 -121
rect -2351 -2109 -2293 -2097
rect -2093 -121 -2035 -109
rect -2093 -2097 -2081 -121
rect -2047 -2097 -2035 -121
rect -2093 -2109 -2035 -2097
rect -1835 -121 -1777 -109
rect -1835 -2097 -1823 -121
rect -1789 -2097 -1777 -121
rect -1835 -2109 -1777 -2097
rect -1577 -121 -1519 -109
rect -1577 -2097 -1565 -121
rect -1531 -2097 -1519 -121
rect -1577 -2109 -1519 -2097
rect -1319 -121 -1261 -109
rect -1319 -2097 -1307 -121
rect -1273 -2097 -1261 -121
rect -1319 -2109 -1261 -2097
rect -1061 -121 -1003 -109
rect -1061 -2097 -1049 -121
rect -1015 -2097 -1003 -121
rect -1061 -2109 -1003 -2097
rect -803 -121 -745 -109
rect -803 -2097 -791 -121
rect -757 -2097 -745 -121
rect -803 -2109 -745 -2097
rect -545 -121 -487 -109
rect -545 -2097 -533 -121
rect -499 -2097 -487 -121
rect -545 -2109 -487 -2097
rect -287 -121 -229 -109
rect -287 -2097 -275 -121
rect -241 -2097 -229 -121
rect -287 -2109 -229 -2097
rect -29 -121 29 -109
rect -29 -2097 -17 -121
rect 17 -2097 29 -121
rect -29 -2109 29 -2097
rect 229 -121 287 -109
rect 229 -2097 241 -121
rect 275 -2097 287 -121
rect 229 -2109 287 -2097
rect 487 -121 545 -109
rect 487 -2097 499 -121
rect 533 -2097 545 -121
rect 487 -2109 545 -2097
rect 745 -121 803 -109
rect 745 -2097 757 -121
rect 791 -2097 803 -121
rect 745 -2109 803 -2097
rect 1003 -121 1061 -109
rect 1003 -2097 1015 -121
rect 1049 -2097 1061 -121
rect 1003 -2109 1061 -2097
rect 1261 -121 1319 -109
rect 1261 -2097 1273 -121
rect 1307 -2097 1319 -121
rect 1261 -2109 1319 -2097
rect 1519 -121 1577 -109
rect 1519 -2097 1531 -121
rect 1565 -2097 1577 -121
rect 1519 -2109 1577 -2097
rect 1777 -121 1835 -109
rect 1777 -2097 1789 -121
rect 1823 -2097 1835 -121
rect 1777 -2109 1835 -2097
rect 2035 -121 2093 -109
rect 2035 -2097 2047 -121
rect 2081 -2097 2093 -121
rect 2035 -2109 2093 -2097
rect 2293 -121 2351 -109
rect 2293 -2097 2305 -121
rect 2339 -2097 2351 -121
rect 2293 -2109 2351 -2097
<< mvndiffc >>
rect -2339 121 -2305 2097
rect -2081 121 -2047 2097
rect -1823 121 -1789 2097
rect -1565 121 -1531 2097
rect -1307 121 -1273 2097
rect -1049 121 -1015 2097
rect -791 121 -757 2097
rect -533 121 -499 2097
rect -275 121 -241 2097
rect -17 121 17 2097
rect 241 121 275 2097
rect 499 121 533 2097
rect 757 121 791 2097
rect 1015 121 1049 2097
rect 1273 121 1307 2097
rect 1531 121 1565 2097
rect 1789 121 1823 2097
rect 2047 121 2081 2097
rect 2305 121 2339 2097
rect -2339 -2097 -2305 -121
rect -2081 -2097 -2047 -121
rect -1823 -2097 -1789 -121
rect -1565 -2097 -1531 -121
rect -1307 -2097 -1273 -121
rect -1049 -2097 -1015 -121
rect -791 -2097 -757 -121
rect -533 -2097 -499 -121
rect -275 -2097 -241 -121
rect -17 -2097 17 -121
rect 241 -2097 275 -121
rect 499 -2097 533 -121
rect 757 -2097 791 -121
rect 1015 -2097 1049 -121
rect 1273 -2097 1307 -121
rect 1531 -2097 1565 -121
rect 1789 -2097 1823 -121
rect 2047 -2097 2081 -121
rect 2305 -2097 2339 -121
<< mvpsubdiff >>
rect -2485 2319 2485 2331
rect -2485 2285 -2377 2319
rect 2377 2285 2485 2319
rect -2485 2273 2485 2285
rect -2485 2223 -2427 2273
rect -2485 -2223 -2473 2223
rect -2439 -2223 -2427 2223
rect 2427 2223 2485 2273
rect -2485 -2273 -2427 -2223
rect 2427 -2223 2439 2223
rect 2473 -2223 2485 2223
rect 2427 -2273 2485 -2223
rect -2485 -2285 2485 -2273
rect -2485 -2319 -2377 -2285
rect 2377 -2319 2485 -2285
rect -2485 -2331 2485 -2319
<< mvpsubdiffcont >>
rect -2377 2285 2377 2319
rect -2473 -2223 -2439 2223
rect 2439 -2223 2473 2223
rect -2377 -2319 2377 -2285
<< poly >>
rect -2293 2181 -2093 2197
rect -2293 2147 -2277 2181
rect -2109 2147 -2093 2181
rect -2293 2109 -2093 2147
rect -2035 2181 -1835 2197
rect -2035 2147 -2019 2181
rect -1851 2147 -1835 2181
rect -2035 2109 -1835 2147
rect -1777 2181 -1577 2197
rect -1777 2147 -1761 2181
rect -1593 2147 -1577 2181
rect -1777 2109 -1577 2147
rect -1519 2181 -1319 2197
rect -1519 2147 -1503 2181
rect -1335 2147 -1319 2181
rect -1519 2109 -1319 2147
rect -1261 2181 -1061 2197
rect -1261 2147 -1245 2181
rect -1077 2147 -1061 2181
rect -1261 2109 -1061 2147
rect -1003 2181 -803 2197
rect -1003 2147 -987 2181
rect -819 2147 -803 2181
rect -1003 2109 -803 2147
rect -745 2181 -545 2197
rect -745 2147 -729 2181
rect -561 2147 -545 2181
rect -745 2109 -545 2147
rect -487 2181 -287 2197
rect -487 2147 -471 2181
rect -303 2147 -287 2181
rect -487 2109 -287 2147
rect -229 2181 -29 2197
rect -229 2147 -213 2181
rect -45 2147 -29 2181
rect -229 2109 -29 2147
rect 29 2181 229 2197
rect 29 2147 45 2181
rect 213 2147 229 2181
rect 29 2109 229 2147
rect 287 2181 487 2197
rect 287 2147 303 2181
rect 471 2147 487 2181
rect 287 2109 487 2147
rect 545 2181 745 2197
rect 545 2147 561 2181
rect 729 2147 745 2181
rect 545 2109 745 2147
rect 803 2181 1003 2197
rect 803 2147 819 2181
rect 987 2147 1003 2181
rect 803 2109 1003 2147
rect 1061 2181 1261 2197
rect 1061 2147 1077 2181
rect 1245 2147 1261 2181
rect 1061 2109 1261 2147
rect 1319 2181 1519 2197
rect 1319 2147 1335 2181
rect 1503 2147 1519 2181
rect 1319 2109 1519 2147
rect 1577 2181 1777 2197
rect 1577 2147 1593 2181
rect 1761 2147 1777 2181
rect 1577 2109 1777 2147
rect 1835 2181 2035 2197
rect 1835 2147 1851 2181
rect 2019 2147 2035 2181
rect 1835 2109 2035 2147
rect 2093 2181 2293 2197
rect 2093 2147 2109 2181
rect 2277 2147 2293 2181
rect 2093 2109 2293 2147
rect -2293 71 -2093 109
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2293 21 -2093 37
rect -2035 71 -1835 109
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 109
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 109
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 109
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 109
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 109
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 109
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 109
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect 2093 71 2293 109
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2093 21 2293 37
rect -2293 -37 -2093 -21
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2293 -109 -2093 -71
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -109 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -109 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -109 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -109 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -109 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -109 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -109 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -109 2035 -71
rect 2093 -37 2293 -21
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2093 -109 2293 -71
rect -2293 -2147 -2093 -2109
rect -2293 -2181 -2277 -2147
rect -2109 -2181 -2093 -2147
rect -2293 -2197 -2093 -2181
rect -2035 -2147 -1835 -2109
rect -2035 -2181 -2019 -2147
rect -1851 -2181 -1835 -2147
rect -2035 -2197 -1835 -2181
rect -1777 -2147 -1577 -2109
rect -1777 -2181 -1761 -2147
rect -1593 -2181 -1577 -2147
rect -1777 -2197 -1577 -2181
rect -1519 -2147 -1319 -2109
rect -1519 -2181 -1503 -2147
rect -1335 -2181 -1319 -2147
rect -1519 -2197 -1319 -2181
rect -1261 -2147 -1061 -2109
rect -1261 -2181 -1245 -2147
rect -1077 -2181 -1061 -2147
rect -1261 -2197 -1061 -2181
rect -1003 -2147 -803 -2109
rect -1003 -2181 -987 -2147
rect -819 -2181 -803 -2147
rect -1003 -2197 -803 -2181
rect -745 -2147 -545 -2109
rect -745 -2181 -729 -2147
rect -561 -2181 -545 -2147
rect -745 -2197 -545 -2181
rect -487 -2147 -287 -2109
rect -487 -2181 -471 -2147
rect -303 -2181 -287 -2147
rect -487 -2197 -287 -2181
rect -229 -2147 -29 -2109
rect -229 -2181 -213 -2147
rect -45 -2181 -29 -2147
rect -229 -2197 -29 -2181
rect 29 -2147 229 -2109
rect 29 -2181 45 -2147
rect 213 -2181 229 -2147
rect 29 -2197 229 -2181
rect 287 -2147 487 -2109
rect 287 -2181 303 -2147
rect 471 -2181 487 -2147
rect 287 -2197 487 -2181
rect 545 -2147 745 -2109
rect 545 -2181 561 -2147
rect 729 -2181 745 -2147
rect 545 -2197 745 -2181
rect 803 -2147 1003 -2109
rect 803 -2181 819 -2147
rect 987 -2181 1003 -2147
rect 803 -2197 1003 -2181
rect 1061 -2147 1261 -2109
rect 1061 -2181 1077 -2147
rect 1245 -2181 1261 -2147
rect 1061 -2197 1261 -2181
rect 1319 -2147 1519 -2109
rect 1319 -2181 1335 -2147
rect 1503 -2181 1519 -2147
rect 1319 -2197 1519 -2181
rect 1577 -2147 1777 -2109
rect 1577 -2181 1593 -2147
rect 1761 -2181 1777 -2147
rect 1577 -2197 1777 -2181
rect 1835 -2147 2035 -2109
rect 1835 -2181 1851 -2147
rect 2019 -2181 2035 -2147
rect 1835 -2197 2035 -2181
rect 2093 -2147 2293 -2109
rect 2093 -2181 2109 -2147
rect 2277 -2181 2293 -2147
rect 2093 -2197 2293 -2181
<< polycont >>
rect -2277 2147 -2109 2181
rect -2019 2147 -1851 2181
rect -1761 2147 -1593 2181
rect -1503 2147 -1335 2181
rect -1245 2147 -1077 2181
rect -987 2147 -819 2181
rect -729 2147 -561 2181
rect -471 2147 -303 2181
rect -213 2147 -45 2181
rect 45 2147 213 2181
rect 303 2147 471 2181
rect 561 2147 729 2181
rect 819 2147 987 2181
rect 1077 2147 1245 2181
rect 1335 2147 1503 2181
rect 1593 2147 1761 2181
rect 1851 2147 2019 2181
rect 2109 2147 2277 2181
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect -2277 -2181 -2109 -2147
rect -2019 -2181 -1851 -2147
rect -1761 -2181 -1593 -2147
rect -1503 -2181 -1335 -2147
rect -1245 -2181 -1077 -2147
rect -987 -2181 -819 -2147
rect -729 -2181 -561 -2147
rect -471 -2181 -303 -2147
rect -213 -2181 -45 -2147
rect 45 -2181 213 -2147
rect 303 -2181 471 -2147
rect 561 -2181 729 -2147
rect 819 -2181 987 -2147
rect 1077 -2181 1245 -2147
rect 1335 -2181 1503 -2147
rect 1593 -2181 1761 -2147
rect 1851 -2181 2019 -2147
rect 2109 -2181 2277 -2147
<< locali >>
rect -2473 2285 -2377 2319
rect 2377 2285 2473 2319
rect -2473 2223 -2439 2285
rect 2439 2223 2473 2285
rect -2293 2147 -2277 2181
rect -2109 2147 -2093 2181
rect -2035 2147 -2019 2181
rect -1851 2147 -1835 2181
rect -1777 2147 -1761 2181
rect -1593 2147 -1577 2181
rect -1519 2147 -1503 2181
rect -1335 2147 -1319 2181
rect -1261 2147 -1245 2181
rect -1077 2147 -1061 2181
rect -1003 2147 -987 2181
rect -819 2147 -803 2181
rect -745 2147 -729 2181
rect -561 2147 -545 2181
rect -487 2147 -471 2181
rect -303 2147 -287 2181
rect -229 2147 -213 2181
rect -45 2147 -29 2181
rect 29 2147 45 2181
rect 213 2147 229 2181
rect 287 2147 303 2181
rect 471 2147 487 2181
rect 545 2147 561 2181
rect 729 2147 745 2181
rect 803 2147 819 2181
rect 987 2147 1003 2181
rect 1061 2147 1077 2181
rect 1245 2147 1261 2181
rect 1319 2147 1335 2181
rect 1503 2147 1519 2181
rect 1577 2147 1593 2181
rect 1761 2147 1777 2181
rect 1835 2147 1851 2181
rect 2019 2147 2035 2181
rect 2093 2147 2109 2181
rect 2277 2147 2293 2181
rect -2339 2097 -2305 2113
rect -2339 105 -2305 121
rect -2081 2097 -2047 2113
rect -2081 105 -2047 121
rect -1823 2097 -1789 2113
rect -1823 105 -1789 121
rect -1565 2097 -1531 2113
rect -1565 105 -1531 121
rect -1307 2097 -1273 2113
rect -1307 105 -1273 121
rect -1049 2097 -1015 2113
rect -1049 105 -1015 121
rect -791 2097 -757 2113
rect -791 105 -757 121
rect -533 2097 -499 2113
rect -533 105 -499 121
rect -275 2097 -241 2113
rect -275 105 -241 121
rect -17 2097 17 2113
rect -17 105 17 121
rect 241 2097 275 2113
rect 241 105 275 121
rect 499 2097 533 2113
rect 499 105 533 121
rect 757 2097 791 2113
rect 757 105 791 121
rect 1015 2097 1049 2113
rect 1015 105 1049 121
rect 1273 2097 1307 2113
rect 1273 105 1307 121
rect 1531 2097 1565 2113
rect 1531 105 1565 121
rect 1789 2097 1823 2113
rect 1789 105 1823 121
rect 2047 2097 2081 2113
rect 2047 105 2081 121
rect 2305 2097 2339 2113
rect 2305 105 2339 121
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 2093 37 2109 71
rect 2277 37 2293 71
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect -2339 -121 -2305 -105
rect -2339 -2113 -2305 -2097
rect -2081 -121 -2047 -105
rect -2081 -2113 -2047 -2097
rect -1823 -121 -1789 -105
rect -1823 -2113 -1789 -2097
rect -1565 -121 -1531 -105
rect -1565 -2113 -1531 -2097
rect -1307 -121 -1273 -105
rect -1307 -2113 -1273 -2097
rect -1049 -121 -1015 -105
rect -1049 -2113 -1015 -2097
rect -791 -121 -757 -105
rect -791 -2113 -757 -2097
rect -533 -121 -499 -105
rect -533 -2113 -499 -2097
rect -275 -121 -241 -105
rect -275 -2113 -241 -2097
rect -17 -121 17 -105
rect -17 -2113 17 -2097
rect 241 -121 275 -105
rect 241 -2113 275 -2097
rect 499 -121 533 -105
rect 499 -2113 533 -2097
rect 757 -121 791 -105
rect 757 -2113 791 -2097
rect 1015 -121 1049 -105
rect 1015 -2113 1049 -2097
rect 1273 -121 1307 -105
rect 1273 -2113 1307 -2097
rect 1531 -121 1565 -105
rect 1531 -2113 1565 -2097
rect 1789 -121 1823 -105
rect 1789 -2113 1823 -2097
rect 2047 -121 2081 -105
rect 2047 -2113 2081 -2097
rect 2305 -121 2339 -105
rect 2305 -2113 2339 -2097
rect -2293 -2181 -2277 -2147
rect -2109 -2181 -2093 -2147
rect -2035 -2181 -2019 -2147
rect -1851 -2181 -1835 -2147
rect -1777 -2181 -1761 -2147
rect -1593 -2181 -1577 -2147
rect -1519 -2181 -1503 -2147
rect -1335 -2181 -1319 -2147
rect -1261 -2181 -1245 -2147
rect -1077 -2181 -1061 -2147
rect -1003 -2181 -987 -2147
rect -819 -2181 -803 -2147
rect -745 -2181 -729 -2147
rect -561 -2181 -545 -2147
rect -487 -2181 -471 -2147
rect -303 -2181 -287 -2147
rect -229 -2181 -213 -2147
rect -45 -2181 -29 -2147
rect 29 -2181 45 -2147
rect 213 -2181 229 -2147
rect 287 -2181 303 -2147
rect 471 -2181 487 -2147
rect 545 -2181 561 -2147
rect 729 -2181 745 -2147
rect 803 -2181 819 -2147
rect 987 -2181 1003 -2147
rect 1061 -2181 1077 -2147
rect 1245 -2181 1261 -2147
rect 1319 -2181 1335 -2147
rect 1503 -2181 1519 -2147
rect 1577 -2181 1593 -2147
rect 1761 -2181 1777 -2147
rect 1835 -2181 1851 -2147
rect 2019 -2181 2035 -2147
rect 2093 -2181 2109 -2147
rect 2277 -2181 2293 -2147
rect -2473 -2285 -2439 -2223
rect 2439 -2285 2473 -2223
rect -2473 -2319 -2377 -2285
rect 2377 -2319 2473 -2285
<< viali >>
rect -2277 2147 -2109 2181
rect -2019 2147 -1851 2181
rect -1761 2147 -1593 2181
rect -1503 2147 -1335 2181
rect -1245 2147 -1077 2181
rect -987 2147 -819 2181
rect -729 2147 -561 2181
rect -471 2147 -303 2181
rect -213 2147 -45 2181
rect 45 2147 213 2181
rect 303 2147 471 2181
rect 561 2147 729 2181
rect 819 2147 987 2181
rect 1077 2147 1245 2181
rect 1335 2147 1503 2181
rect 1593 2147 1761 2181
rect 1851 2147 2019 2181
rect 2109 2147 2277 2181
rect -2339 121 -2305 2097
rect -2081 121 -2047 2097
rect -1823 121 -1789 2097
rect -1565 121 -1531 2097
rect -1307 121 -1273 2097
rect -1049 121 -1015 2097
rect -791 121 -757 2097
rect -533 121 -499 2097
rect -275 121 -241 2097
rect -17 121 17 2097
rect 241 121 275 2097
rect 499 121 533 2097
rect 757 121 791 2097
rect 1015 121 1049 2097
rect 1273 121 1307 2097
rect 1531 121 1565 2097
rect 1789 121 1823 2097
rect 2047 121 2081 2097
rect 2305 121 2339 2097
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect -2339 -2097 -2305 -121
rect -2081 -2097 -2047 -121
rect -1823 -2097 -1789 -121
rect -1565 -2097 -1531 -121
rect -1307 -2097 -1273 -121
rect -1049 -2097 -1015 -121
rect -791 -2097 -757 -121
rect -533 -2097 -499 -121
rect -275 -2097 -241 -121
rect -17 -2097 17 -121
rect 241 -2097 275 -121
rect 499 -2097 533 -121
rect 757 -2097 791 -121
rect 1015 -2097 1049 -121
rect 1273 -2097 1307 -121
rect 1531 -2097 1565 -121
rect 1789 -2097 1823 -121
rect 2047 -2097 2081 -121
rect 2305 -2097 2339 -121
rect -2277 -2181 -2109 -2147
rect -2019 -2181 -1851 -2147
rect -1761 -2181 -1593 -2147
rect -1503 -2181 -1335 -2147
rect -1245 -2181 -1077 -2147
rect -987 -2181 -819 -2147
rect -729 -2181 -561 -2147
rect -471 -2181 -303 -2147
rect -213 -2181 -45 -2147
rect 45 -2181 213 -2147
rect 303 -2181 471 -2147
rect 561 -2181 729 -2147
rect 819 -2181 987 -2147
rect 1077 -2181 1245 -2147
rect 1335 -2181 1503 -2147
rect 1593 -2181 1761 -2147
rect 1851 -2181 2019 -2147
rect 2109 -2181 2277 -2147
<< metal1 >>
rect -2289 2181 -2097 2187
rect -2289 2147 -2277 2181
rect -2109 2147 -2097 2181
rect -2289 2141 -2097 2147
rect -2031 2181 -1839 2187
rect -2031 2147 -2019 2181
rect -1851 2147 -1839 2181
rect -2031 2141 -1839 2147
rect -1773 2181 -1581 2187
rect -1773 2147 -1761 2181
rect -1593 2147 -1581 2181
rect -1773 2141 -1581 2147
rect -1515 2181 -1323 2187
rect -1515 2147 -1503 2181
rect -1335 2147 -1323 2181
rect -1515 2141 -1323 2147
rect -1257 2181 -1065 2187
rect -1257 2147 -1245 2181
rect -1077 2147 -1065 2181
rect -1257 2141 -1065 2147
rect -999 2181 -807 2187
rect -999 2147 -987 2181
rect -819 2147 -807 2181
rect -999 2141 -807 2147
rect -741 2181 -549 2187
rect -741 2147 -729 2181
rect -561 2147 -549 2181
rect -741 2141 -549 2147
rect -483 2181 -291 2187
rect -483 2147 -471 2181
rect -303 2147 -291 2181
rect -483 2141 -291 2147
rect -225 2181 -33 2187
rect -225 2147 -213 2181
rect -45 2147 -33 2181
rect -225 2141 -33 2147
rect 33 2181 225 2187
rect 33 2147 45 2181
rect 213 2147 225 2181
rect 33 2141 225 2147
rect 291 2181 483 2187
rect 291 2147 303 2181
rect 471 2147 483 2181
rect 291 2141 483 2147
rect 549 2181 741 2187
rect 549 2147 561 2181
rect 729 2147 741 2181
rect 549 2141 741 2147
rect 807 2181 999 2187
rect 807 2147 819 2181
rect 987 2147 999 2181
rect 807 2141 999 2147
rect 1065 2181 1257 2187
rect 1065 2147 1077 2181
rect 1245 2147 1257 2181
rect 1065 2141 1257 2147
rect 1323 2181 1515 2187
rect 1323 2147 1335 2181
rect 1503 2147 1515 2181
rect 1323 2141 1515 2147
rect 1581 2181 1773 2187
rect 1581 2147 1593 2181
rect 1761 2147 1773 2181
rect 1581 2141 1773 2147
rect 1839 2181 2031 2187
rect 1839 2147 1851 2181
rect 2019 2147 2031 2181
rect 1839 2141 2031 2147
rect 2097 2181 2289 2187
rect 2097 2147 2109 2181
rect 2277 2147 2289 2181
rect 2097 2141 2289 2147
rect -2345 2097 -2299 2109
rect -2345 121 -2339 2097
rect -2305 121 -2299 2097
rect -2345 109 -2299 121
rect -2087 2097 -2041 2109
rect -2087 121 -2081 2097
rect -2047 121 -2041 2097
rect -2087 109 -2041 121
rect -1829 2097 -1783 2109
rect -1829 121 -1823 2097
rect -1789 121 -1783 2097
rect -1829 109 -1783 121
rect -1571 2097 -1525 2109
rect -1571 121 -1565 2097
rect -1531 121 -1525 2097
rect -1571 109 -1525 121
rect -1313 2097 -1267 2109
rect -1313 121 -1307 2097
rect -1273 121 -1267 2097
rect -1313 109 -1267 121
rect -1055 2097 -1009 2109
rect -1055 121 -1049 2097
rect -1015 121 -1009 2097
rect -1055 109 -1009 121
rect -797 2097 -751 2109
rect -797 121 -791 2097
rect -757 121 -751 2097
rect -797 109 -751 121
rect -539 2097 -493 2109
rect -539 121 -533 2097
rect -499 121 -493 2097
rect -539 109 -493 121
rect -281 2097 -235 2109
rect -281 121 -275 2097
rect -241 121 -235 2097
rect -281 109 -235 121
rect -23 2097 23 2109
rect -23 121 -17 2097
rect 17 121 23 2097
rect -23 109 23 121
rect 235 2097 281 2109
rect 235 121 241 2097
rect 275 121 281 2097
rect 235 109 281 121
rect 493 2097 539 2109
rect 493 121 499 2097
rect 533 121 539 2097
rect 493 109 539 121
rect 751 2097 797 2109
rect 751 121 757 2097
rect 791 121 797 2097
rect 751 109 797 121
rect 1009 2097 1055 2109
rect 1009 121 1015 2097
rect 1049 121 1055 2097
rect 1009 109 1055 121
rect 1267 2097 1313 2109
rect 1267 121 1273 2097
rect 1307 121 1313 2097
rect 1267 109 1313 121
rect 1525 2097 1571 2109
rect 1525 121 1531 2097
rect 1565 121 1571 2097
rect 1525 109 1571 121
rect 1783 2097 1829 2109
rect 1783 121 1789 2097
rect 1823 121 1829 2097
rect 1783 109 1829 121
rect 2041 2097 2087 2109
rect 2041 121 2047 2097
rect 2081 121 2087 2097
rect 2041 109 2087 121
rect 2299 2097 2345 2109
rect 2299 121 2305 2097
rect 2339 121 2345 2097
rect 2299 109 2345 121
rect -2289 71 -2097 77
rect -2289 37 -2277 71
rect -2109 37 -2097 71
rect -2289 31 -2097 37
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect 2097 71 2289 77
rect 2097 37 2109 71
rect 2277 37 2289 71
rect 2097 31 2289 37
rect -2289 -37 -2097 -31
rect -2289 -71 -2277 -37
rect -2109 -71 -2097 -37
rect -2289 -77 -2097 -71
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect 2097 -37 2289 -31
rect 2097 -71 2109 -37
rect 2277 -71 2289 -37
rect 2097 -77 2289 -71
rect -2345 -121 -2299 -109
rect -2345 -2097 -2339 -121
rect -2305 -2097 -2299 -121
rect -2345 -2109 -2299 -2097
rect -2087 -121 -2041 -109
rect -2087 -2097 -2081 -121
rect -2047 -2097 -2041 -121
rect -2087 -2109 -2041 -2097
rect -1829 -121 -1783 -109
rect -1829 -2097 -1823 -121
rect -1789 -2097 -1783 -121
rect -1829 -2109 -1783 -2097
rect -1571 -121 -1525 -109
rect -1571 -2097 -1565 -121
rect -1531 -2097 -1525 -121
rect -1571 -2109 -1525 -2097
rect -1313 -121 -1267 -109
rect -1313 -2097 -1307 -121
rect -1273 -2097 -1267 -121
rect -1313 -2109 -1267 -2097
rect -1055 -121 -1009 -109
rect -1055 -2097 -1049 -121
rect -1015 -2097 -1009 -121
rect -1055 -2109 -1009 -2097
rect -797 -121 -751 -109
rect -797 -2097 -791 -121
rect -757 -2097 -751 -121
rect -797 -2109 -751 -2097
rect -539 -121 -493 -109
rect -539 -2097 -533 -121
rect -499 -2097 -493 -121
rect -539 -2109 -493 -2097
rect -281 -121 -235 -109
rect -281 -2097 -275 -121
rect -241 -2097 -235 -121
rect -281 -2109 -235 -2097
rect -23 -121 23 -109
rect -23 -2097 -17 -121
rect 17 -2097 23 -121
rect -23 -2109 23 -2097
rect 235 -121 281 -109
rect 235 -2097 241 -121
rect 275 -2097 281 -121
rect 235 -2109 281 -2097
rect 493 -121 539 -109
rect 493 -2097 499 -121
rect 533 -2097 539 -121
rect 493 -2109 539 -2097
rect 751 -121 797 -109
rect 751 -2097 757 -121
rect 791 -2097 797 -121
rect 751 -2109 797 -2097
rect 1009 -121 1055 -109
rect 1009 -2097 1015 -121
rect 1049 -2097 1055 -121
rect 1009 -2109 1055 -2097
rect 1267 -121 1313 -109
rect 1267 -2097 1273 -121
rect 1307 -2097 1313 -121
rect 1267 -2109 1313 -2097
rect 1525 -121 1571 -109
rect 1525 -2097 1531 -121
rect 1565 -2097 1571 -121
rect 1525 -2109 1571 -2097
rect 1783 -121 1829 -109
rect 1783 -2097 1789 -121
rect 1823 -2097 1829 -121
rect 1783 -2109 1829 -2097
rect 2041 -121 2087 -109
rect 2041 -2097 2047 -121
rect 2081 -2097 2087 -121
rect 2041 -2109 2087 -2097
rect 2299 -121 2345 -109
rect 2299 -2097 2305 -121
rect 2339 -2097 2345 -121
rect 2299 -2109 2345 -2097
rect -2289 -2147 -2097 -2141
rect -2289 -2181 -2277 -2147
rect -2109 -2181 -2097 -2147
rect -2289 -2187 -2097 -2181
rect -2031 -2147 -1839 -2141
rect -2031 -2181 -2019 -2147
rect -1851 -2181 -1839 -2147
rect -2031 -2187 -1839 -2181
rect -1773 -2147 -1581 -2141
rect -1773 -2181 -1761 -2147
rect -1593 -2181 -1581 -2147
rect -1773 -2187 -1581 -2181
rect -1515 -2147 -1323 -2141
rect -1515 -2181 -1503 -2147
rect -1335 -2181 -1323 -2147
rect -1515 -2187 -1323 -2181
rect -1257 -2147 -1065 -2141
rect -1257 -2181 -1245 -2147
rect -1077 -2181 -1065 -2147
rect -1257 -2187 -1065 -2181
rect -999 -2147 -807 -2141
rect -999 -2181 -987 -2147
rect -819 -2181 -807 -2147
rect -999 -2187 -807 -2181
rect -741 -2147 -549 -2141
rect -741 -2181 -729 -2147
rect -561 -2181 -549 -2147
rect -741 -2187 -549 -2181
rect -483 -2147 -291 -2141
rect -483 -2181 -471 -2147
rect -303 -2181 -291 -2147
rect -483 -2187 -291 -2181
rect -225 -2147 -33 -2141
rect -225 -2181 -213 -2147
rect -45 -2181 -33 -2147
rect -225 -2187 -33 -2181
rect 33 -2147 225 -2141
rect 33 -2181 45 -2147
rect 213 -2181 225 -2147
rect 33 -2187 225 -2181
rect 291 -2147 483 -2141
rect 291 -2181 303 -2147
rect 471 -2181 483 -2147
rect 291 -2187 483 -2181
rect 549 -2147 741 -2141
rect 549 -2181 561 -2147
rect 729 -2181 741 -2147
rect 549 -2187 741 -2181
rect 807 -2147 999 -2141
rect 807 -2181 819 -2147
rect 987 -2181 999 -2147
rect 807 -2187 999 -2181
rect 1065 -2147 1257 -2141
rect 1065 -2181 1077 -2147
rect 1245 -2181 1257 -2147
rect 1065 -2187 1257 -2181
rect 1323 -2147 1515 -2141
rect 1323 -2181 1335 -2147
rect 1503 -2181 1515 -2147
rect 1323 -2187 1515 -2181
rect 1581 -2147 1773 -2141
rect 1581 -2181 1593 -2147
rect 1761 -2181 1773 -2147
rect 1581 -2187 1773 -2181
rect 1839 -2147 2031 -2141
rect 1839 -2181 1851 -2147
rect 2019 -2181 2031 -2147
rect 1839 -2187 2031 -2181
rect 2097 -2147 2289 -2141
rect 2097 -2181 2109 -2147
rect 2277 -2181 2289 -2147
rect 2097 -2187 2289 -2181
<< properties >>
string FIXED_BBOX -2456 -2302 2456 2302
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10 l 1 m 2 nf 18 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713406689
<< metal3 >>
rect -8916 8012 -6144 8040
rect -8916 5588 -6228 8012
rect -6164 5588 -6144 8012
rect -8916 5560 -6144 5588
rect -5904 8012 -3132 8040
rect -5904 5588 -3216 8012
rect -3152 5588 -3132 8012
rect -5904 5560 -3132 5588
rect -2892 8012 -120 8040
rect -2892 5588 -204 8012
rect -140 5588 -120 8012
rect -2892 5560 -120 5588
rect 120 8012 2892 8040
rect 120 5588 2808 8012
rect 2872 5588 2892 8012
rect 120 5560 2892 5588
rect 3132 8012 5904 8040
rect 3132 5588 5820 8012
rect 5884 5588 5904 8012
rect 3132 5560 5904 5588
rect 6144 8012 8916 8040
rect 6144 5588 8832 8012
rect 8896 5588 8916 8012
rect 6144 5560 8916 5588
rect -8916 5292 -6144 5320
rect -8916 2868 -6228 5292
rect -6164 2868 -6144 5292
rect -8916 2840 -6144 2868
rect -5904 5292 -3132 5320
rect -5904 2868 -3216 5292
rect -3152 2868 -3132 5292
rect -5904 2840 -3132 2868
rect -2892 5292 -120 5320
rect -2892 2868 -204 5292
rect -140 2868 -120 5292
rect -2892 2840 -120 2868
rect 120 5292 2892 5320
rect 120 2868 2808 5292
rect 2872 2868 2892 5292
rect 120 2840 2892 2868
rect 3132 5292 5904 5320
rect 3132 2868 5820 5292
rect 5884 2868 5904 5292
rect 3132 2840 5904 2868
rect 6144 5292 8916 5320
rect 6144 2868 8832 5292
rect 8896 2868 8916 5292
rect 6144 2840 8916 2868
rect -8916 2572 -6144 2600
rect -8916 148 -6228 2572
rect -6164 148 -6144 2572
rect -8916 120 -6144 148
rect -5904 2572 -3132 2600
rect -5904 148 -3216 2572
rect -3152 148 -3132 2572
rect -5904 120 -3132 148
rect -2892 2572 -120 2600
rect -2892 148 -204 2572
rect -140 148 -120 2572
rect -2892 120 -120 148
rect 120 2572 2892 2600
rect 120 148 2808 2572
rect 2872 148 2892 2572
rect 120 120 2892 148
rect 3132 2572 5904 2600
rect 3132 148 5820 2572
rect 5884 148 5904 2572
rect 3132 120 5904 148
rect 6144 2572 8916 2600
rect 6144 148 8832 2572
rect 8896 148 8916 2572
rect 6144 120 8916 148
rect -8916 -148 -6144 -120
rect -8916 -2572 -6228 -148
rect -6164 -2572 -6144 -148
rect -8916 -2600 -6144 -2572
rect -5904 -148 -3132 -120
rect -5904 -2572 -3216 -148
rect -3152 -2572 -3132 -148
rect -5904 -2600 -3132 -2572
rect -2892 -148 -120 -120
rect -2892 -2572 -204 -148
rect -140 -2572 -120 -148
rect -2892 -2600 -120 -2572
rect 120 -148 2892 -120
rect 120 -2572 2808 -148
rect 2872 -2572 2892 -148
rect 120 -2600 2892 -2572
rect 3132 -148 5904 -120
rect 3132 -2572 5820 -148
rect 5884 -2572 5904 -148
rect 3132 -2600 5904 -2572
rect 6144 -148 8916 -120
rect 6144 -2572 8832 -148
rect 8896 -2572 8916 -148
rect 6144 -2600 8916 -2572
rect -8916 -2868 -6144 -2840
rect -8916 -5292 -6228 -2868
rect -6164 -5292 -6144 -2868
rect -8916 -5320 -6144 -5292
rect -5904 -2868 -3132 -2840
rect -5904 -5292 -3216 -2868
rect -3152 -5292 -3132 -2868
rect -5904 -5320 -3132 -5292
rect -2892 -2868 -120 -2840
rect -2892 -5292 -204 -2868
rect -140 -5292 -120 -2868
rect -2892 -5320 -120 -5292
rect 120 -2868 2892 -2840
rect 120 -5292 2808 -2868
rect 2872 -5292 2892 -2868
rect 120 -5320 2892 -5292
rect 3132 -2868 5904 -2840
rect 3132 -5292 5820 -2868
rect 5884 -5292 5904 -2868
rect 3132 -5320 5904 -5292
rect 6144 -2868 8916 -2840
rect 6144 -5292 8832 -2868
rect 8896 -5292 8916 -2868
rect 6144 -5320 8916 -5292
rect -8916 -5588 -6144 -5560
rect -8916 -8012 -6228 -5588
rect -6164 -8012 -6144 -5588
rect -8916 -8040 -6144 -8012
rect -5904 -5588 -3132 -5560
rect -5904 -8012 -3216 -5588
rect -3152 -8012 -3132 -5588
rect -5904 -8040 -3132 -8012
rect -2892 -5588 -120 -5560
rect -2892 -8012 -204 -5588
rect -140 -8012 -120 -5588
rect -2892 -8040 -120 -8012
rect 120 -5588 2892 -5560
rect 120 -8012 2808 -5588
rect 2872 -8012 2892 -5588
rect 120 -8040 2892 -8012
rect 3132 -5588 5904 -5560
rect 3132 -8012 5820 -5588
rect 5884 -8012 5904 -5588
rect 3132 -8040 5904 -8012
rect 6144 -5588 8916 -5560
rect 6144 -8012 8832 -5588
rect 8896 -8012 8916 -5588
rect 6144 -8040 8916 -8012
<< via3 >>
rect -6228 5588 -6164 8012
rect -3216 5588 -3152 8012
rect -204 5588 -140 8012
rect 2808 5588 2872 8012
rect 5820 5588 5884 8012
rect 8832 5588 8896 8012
rect -6228 2868 -6164 5292
rect -3216 2868 -3152 5292
rect -204 2868 -140 5292
rect 2808 2868 2872 5292
rect 5820 2868 5884 5292
rect 8832 2868 8896 5292
rect -6228 148 -6164 2572
rect -3216 148 -3152 2572
rect -204 148 -140 2572
rect 2808 148 2872 2572
rect 5820 148 5884 2572
rect 8832 148 8896 2572
rect -6228 -2572 -6164 -148
rect -3216 -2572 -3152 -148
rect -204 -2572 -140 -148
rect 2808 -2572 2872 -148
rect 5820 -2572 5884 -148
rect 8832 -2572 8896 -148
rect -6228 -5292 -6164 -2868
rect -3216 -5292 -3152 -2868
rect -204 -5292 -140 -2868
rect 2808 -5292 2872 -2868
rect 5820 -5292 5884 -2868
rect 8832 -5292 8896 -2868
rect -6228 -8012 -6164 -5588
rect -3216 -8012 -3152 -5588
rect -204 -8012 -140 -5588
rect 2808 -8012 2872 -5588
rect 5820 -8012 5884 -5588
rect 8832 -8012 8896 -5588
<< mimcap >>
rect -8876 7960 -6476 8000
rect -8876 5640 -8836 7960
rect -6516 5640 -6476 7960
rect -8876 5600 -6476 5640
rect -5864 7960 -3464 8000
rect -5864 5640 -5824 7960
rect -3504 5640 -3464 7960
rect -5864 5600 -3464 5640
rect -2852 7960 -452 8000
rect -2852 5640 -2812 7960
rect -492 5640 -452 7960
rect -2852 5600 -452 5640
rect 160 7960 2560 8000
rect 160 5640 200 7960
rect 2520 5640 2560 7960
rect 160 5600 2560 5640
rect 3172 7960 5572 8000
rect 3172 5640 3212 7960
rect 5532 5640 5572 7960
rect 3172 5600 5572 5640
rect 6184 7960 8584 8000
rect 6184 5640 6224 7960
rect 8544 5640 8584 7960
rect 6184 5600 8584 5640
rect -8876 5240 -6476 5280
rect -8876 2920 -8836 5240
rect -6516 2920 -6476 5240
rect -8876 2880 -6476 2920
rect -5864 5240 -3464 5280
rect -5864 2920 -5824 5240
rect -3504 2920 -3464 5240
rect -5864 2880 -3464 2920
rect -2852 5240 -452 5280
rect -2852 2920 -2812 5240
rect -492 2920 -452 5240
rect -2852 2880 -452 2920
rect 160 5240 2560 5280
rect 160 2920 200 5240
rect 2520 2920 2560 5240
rect 160 2880 2560 2920
rect 3172 5240 5572 5280
rect 3172 2920 3212 5240
rect 5532 2920 5572 5240
rect 3172 2880 5572 2920
rect 6184 5240 8584 5280
rect 6184 2920 6224 5240
rect 8544 2920 8584 5240
rect 6184 2880 8584 2920
rect -8876 2520 -6476 2560
rect -8876 200 -8836 2520
rect -6516 200 -6476 2520
rect -8876 160 -6476 200
rect -5864 2520 -3464 2560
rect -5864 200 -5824 2520
rect -3504 200 -3464 2520
rect -5864 160 -3464 200
rect -2852 2520 -452 2560
rect -2852 200 -2812 2520
rect -492 200 -452 2520
rect -2852 160 -452 200
rect 160 2520 2560 2560
rect 160 200 200 2520
rect 2520 200 2560 2520
rect 160 160 2560 200
rect 3172 2520 5572 2560
rect 3172 200 3212 2520
rect 5532 200 5572 2520
rect 3172 160 5572 200
rect 6184 2520 8584 2560
rect 6184 200 6224 2520
rect 8544 200 8584 2520
rect 6184 160 8584 200
rect -8876 -200 -6476 -160
rect -8876 -2520 -8836 -200
rect -6516 -2520 -6476 -200
rect -8876 -2560 -6476 -2520
rect -5864 -200 -3464 -160
rect -5864 -2520 -5824 -200
rect -3504 -2520 -3464 -200
rect -5864 -2560 -3464 -2520
rect -2852 -200 -452 -160
rect -2852 -2520 -2812 -200
rect -492 -2520 -452 -200
rect -2852 -2560 -452 -2520
rect 160 -200 2560 -160
rect 160 -2520 200 -200
rect 2520 -2520 2560 -200
rect 160 -2560 2560 -2520
rect 3172 -200 5572 -160
rect 3172 -2520 3212 -200
rect 5532 -2520 5572 -200
rect 3172 -2560 5572 -2520
rect 6184 -200 8584 -160
rect 6184 -2520 6224 -200
rect 8544 -2520 8584 -200
rect 6184 -2560 8584 -2520
rect -8876 -2920 -6476 -2880
rect -8876 -5240 -8836 -2920
rect -6516 -5240 -6476 -2920
rect -8876 -5280 -6476 -5240
rect -5864 -2920 -3464 -2880
rect -5864 -5240 -5824 -2920
rect -3504 -5240 -3464 -2920
rect -5864 -5280 -3464 -5240
rect -2852 -2920 -452 -2880
rect -2852 -5240 -2812 -2920
rect -492 -5240 -452 -2920
rect -2852 -5280 -452 -5240
rect 160 -2920 2560 -2880
rect 160 -5240 200 -2920
rect 2520 -5240 2560 -2920
rect 160 -5280 2560 -5240
rect 3172 -2920 5572 -2880
rect 3172 -5240 3212 -2920
rect 5532 -5240 5572 -2920
rect 3172 -5280 5572 -5240
rect 6184 -2920 8584 -2880
rect 6184 -5240 6224 -2920
rect 8544 -5240 8584 -2920
rect 6184 -5280 8584 -5240
rect -8876 -5640 -6476 -5600
rect -8876 -7960 -8836 -5640
rect -6516 -7960 -6476 -5640
rect -8876 -8000 -6476 -7960
rect -5864 -5640 -3464 -5600
rect -5864 -7960 -5824 -5640
rect -3504 -7960 -3464 -5640
rect -5864 -8000 -3464 -7960
rect -2852 -5640 -452 -5600
rect -2852 -7960 -2812 -5640
rect -492 -7960 -452 -5640
rect -2852 -8000 -452 -7960
rect 160 -5640 2560 -5600
rect 160 -7960 200 -5640
rect 2520 -7960 2560 -5640
rect 160 -8000 2560 -7960
rect 3172 -5640 5572 -5600
rect 3172 -7960 3212 -5640
rect 5532 -7960 5572 -5640
rect 3172 -8000 5572 -7960
rect 6184 -5640 8584 -5600
rect 6184 -7960 6224 -5640
rect 8544 -7960 8584 -5640
rect 6184 -8000 8584 -7960
<< mimcapcontact >>
rect -8836 5640 -6516 7960
rect -5824 5640 -3504 7960
rect -2812 5640 -492 7960
rect 200 5640 2520 7960
rect 3212 5640 5532 7960
rect 6224 5640 8544 7960
rect -8836 2920 -6516 5240
rect -5824 2920 -3504 5240
rect -2812 2920 -492 5240
rect 200 2920 2520 5240
rect 3212 2920 5532 5240
rect 6224 2920 8544 5240
rect -8836 200 -6516 2520
rect -5824 200 -3504 2520
rect -2812 200 -492 2520
rect 200 200 2520 2520
rect 3212 200 5532 2520
rect 6224 200 8544 2520
rect -8836 -2520 -6516 -200
rect -5824 -2520 -3504 -200
rect -2812 -2520 -492 -200
rect 200 -2520 2520 -200
rect 3212 -2520 5532 -200
rect 6224 -2520 8544 -200
rect -8836 -5240 -6516 -2920
rect -5824 -5240 -3504 -2920
rect -2812 -5240 -492 -2920
rect 200 -5240 2520 -2920
rect 3212 -5240 5532 -2920
rect 6224 -5240 8544 -2920
rect -8836 -7960 -6516 -5640
rect -5824 -7960 -3504 -5640
rect -2812 -7960 -492 -5640
rect 200 -7960 2520 -5640
rect 3212 -7960 5532 -5640
rect 6224 -7960 8544 -5640
<< metal4 >>
rect -6244 8012 -6148 8028
rect -8837 7960 -6515 7961
rect -8837 5640 -8836 7960
rect -6516 5640 -6515 7960
rect -8837 5639 -6515 5640
rect -6244 5588 -6228 8012
rect -6164 5588 -6148 8012
rect -3232 8012 -3136 8028
rect -5825 7960 -3503 7961
rect -5825 5640 -5824 7960
rect -3504 5640 -3503 7960
rect -5825 5639 -3503 5640
rect -6244 5572 -6148 5588
rect -3232 5588 -3216 8012
rect -3152 5588 -3136 8012
rect -220 8012 -124 8028
rect -2813 7960 -491 7961
rect -2813 5640 -2812 7960
rect -492 5640 -491 7960
rect -2813 5639 -491 5640
rect -3232 5572 -3136 5588
rect -220 5588 -204 8012
rect -140 5588 -124 8012
rect 2792 8012 2888 8028
rect 199 7960 2521 7961
rect 199 5640 200 7960
rect 2520 5640 2521 7960
rect 199 5639 2521 5640
rect -220 5572 -124 5588
rect 2792 5588 2808 8012
rect 2872 5588 2888 8012
rect 5804 8012 5900 8028
rect 3211 7960 5533 7961
rect 3211 5640 3212 7960
rect 5532 5640 5533 7960
rect 3211 5639 5533 5640
rect 2792 5572 2888 5588
rect 5804 5588 5820 8012
rect 5884 5588 5900 8012
rect 8816 8012 8912 8028
rect 6223 7960 8545 7961
rect 6223 5640 6224 7960
rect 8544 5640 8545 7960
rect 6223 5639 8545 5640
rect 5804 5572 5900 5588
rect 8816 5588 8832 8012
rect 8896 5588 8912 8012
rect 8816 5572 8912 5588
rect -6244 5292 -6148 5308
rect -8837 5240 -6515 5241
rect -8837 2920 -8836 5240
rect -6516 2920 -6515 5240
rect -8837 2919 -6515 2920
rect -6244 2868 -6228 5292
rect -6164 2868 -6148 5292
rect -3232 5292 -3136 5308
rect -5825 5240 -3503 5241
rect -5825 2920 -5824 5240
rect -3504 2920 -3503 5240
rect -5825 2919 -3503 2920
rect -6244 2852 -6148 2868
rect -3232 2868 -3216 5292
rect -3152 2868 -3136 5292
rect -220 5292 -124 5308
rect -2813 5240 -491 5241
rect -2813 2920 -2812 5240
rect -492 2920 -491 5240
rect -2813 2919 -491 2920
rect -3232 2852 -3136 2868
rect -220 2868 -204 5292
rect -140 2868 -124 5292
rect 2792 5292 2888 5308
rect 199 5240 2521 5241
rect 199 2920 200 5240
rect 2520 2920 2521 5240
rect 199 2919 2521 2920
rect -220 2852 -124 2868
rect 2792 2868 2808 5292
rect 2872 2868 2888 5292
rect 5804 5292 5900 5308
rect 3211 5240 5533 5241
rect 3211 2920 3212 5240
rect 5532 2920 5533 5240
rect 3211 2919 5533 2920
rect 2792 2852 2888 2868
rect 5804 2868 5820 5292
rect 5884 2868 5900 5292
rect 8816 5292 8912 5308
rect 6223 5240 8545 5241
rect 6223 2920 6224 5240
rect 8544 2920 8545 5240
rect 6223 2919 8545 2920
rect 5804 2852 5900 2868
rect 8816 2868 8832 5292
rect 8896 2868 8912 5292
rect 8816 2852 8912 2868
rect -6244 2572 -6148 2588
rect -8837 2520 -6515 2521
rect -8837 200 -8836 2520
rect -6516 200 -6515 2520
rect -8837 199 -6515 200
rect -6244 148 -6228 2572
rect -6164 148 -6148 2572
rect -3232 2572 -3136 2588
rect -5825 2520 -3503 2521
rect -5825 200 -5824 2520
rect -3504 200 -3503 2520
rect -5825 199 -3503 200
rect -6244 132 -6148 148
rect -3232 148 -3216 2572
rect -3152 148 -3136 2572
rect -220 2572 -124 2588
rect -2813 2520 -491 2521
rect -2813 200 -2812 2520
rect -492 200 -491 2520
rect -2813 199 -491 200
rect -3232 132 -3136 148
rect -220 148 -204 2572
rect -140 148 -124 2572
rect 2792 2572 2888 2588
rect 199 2520 2521 2521
rect 199 200 200 2520
rect 2520 200 2521 2520
rect 199 199 2521 200
rect -220 132 -124 148
rect 2792 148 2808 2572
rect 2872 148 2888 2572
rect 5804 2572 5900 2588
rect 3211 2520 5533 2521
rect 3211 200 3212 2520
rect 5532 200 5533 2520
rect 3211 199 5533 200
rect 2792 132 2888 148
rect 5804 148 5820 2572
rect 5884 148 5900 2572
rect 8816 2572 8912 2588
rect 6223 2520 8545 2521
rect 6223 200 6224 2520
rect 8544 200 8545 2520
rect 6223 199 8545 200
rect 5804 132 5900 148
rect 8816 148 8832 2572
rect 8896 148 8912 2572
rect 8816 132 8912 148
rect -6244 -148 -6148 -132
rect -8837 -200 -6515 -199
rect -8837 -2520 -8836 -200
rect -6516 -2520 -6515 -200
rect -8837 -2521 -6515 -2520
rect -6244 -2572 -6228 -148
rect -6164 -2572 -6148 -148
rect -3232 -148 -3136 -132
rect -5825 -200 -3503 -199
rect -5825 -2520 -5824 -200
rect -3504 -2520 -3503 -200
rect -5825 -2521 -3503 -2520
rect -6244 -2588 -6148 -2572
rect -3232 -2572 -3216 -148
rect -3152 -2572 -3136 -148
rect -220 -148 -124 -132
rect -2813 -200 -491 -199
rect -2813 -2520 -2812 -200
rect -492 -2520 -491 -200
rect -2813 -2521 -491 -2520
rect -3232 -2588 -3136 -2572
rect -220 -2572 -204 -148
rect -140 -2572 -124 -148
rect 2792 -148 2888 -132
rect 199 -200 2521 -199
rect 199 -2520 200 -200
rect 2520 -2520 2521 -200
rect 199 -2521 2521 -2520
rect -220 -2588 -124 -2572
rect 2792 -2572 2808 -148
rect 2872 -2572 2888 -148
rect 5804 -148 5900 -132
rect 3211 -200 5533 -199
rect 3211 -2520 3212 -200
rect 5532 -2520 5533 -200
rect 3211 -2521 5533 -2520
rect 2792 -2588 2888 -2572
rect 5804 -2572 5820 -148
rect 5884 -2572 5900 -148
rect 8816 -148 8912 -132
rect 6223 -200 8545 -199
rect 6223 -2520 6224 -200
rect 8544 -2520 8545 -200
rect 6223 -2521 8545 -2520
rect 5804 -2588 5900 -2572
rect 8816 -2572 8832 -148
rect 8896 -2572 8912 -148
rect 8816 -2588 8912 -2572
rect -6244 -2868 -6148 -2852
rect -8837 -2920 -6515 -2919
rect -8837 -5240 -8836 -2920
rect -6516 -5240 -6515 -2920
rect -8837 -5241 -6515 -5240
rect -6244 -5292 -6228 -2868
rect -6164 -5292 -6148 -2868
rect -3232 -2868 -3136 -2852
rect -5825 -2920 -3503 -2919
rect -5825 -5240 -5824 -2920
rect -3504 -5240 -3503 -2920
rect -5825 -5241 -3503 -5240
rect -6244 -5308 -6148 -5292
rect -3232 -5292 -3216 -2868
rect -3152 -5292 -3136 -2868
rect -220 -2868 -124 -2852
rect -2813 -2920 -491 -2919
rect -2813 -5240 -2812 -2920
rect -492 -5240 -491 -2920
rect -2813 -5241 -491 -5240
rect -3232 -5308 -3136 -5292
rect -220 -5292 -204 -2868
rect -140 -5292 -124 -2868
rect 2792 -2868 2888 -2852
rect 199 -2920 2521 -2919
rect 199 -5240 200 -2920
rect 2520 -5240 2521 -2920
rect 199 -5241 2521 -5240
rect -220 -5308 -124 -5292
rect 2792 -5292 2808 -2868
rect 2872 -5292 2888 -2868
rect 5804 -2868 5900 -2852
rect 3211 -2920 5533 -2919
rect 3211 -5240 3212 -2920
rect 5532 -5240 5533 -2920
rect 3211 -5241 5533 -5240
rect 2792 -5308 2888 -5292
rect 5804 -5292 5820 -2868
rect 5884 -5292 5900 -2868
rect 8816 -2868 8912 -2852
rect 6223 -2920 8545 -2919
rect 6223 -5240 6224 -2920
rect 8544 -5240 8545 -2920
rect 6223 -5241 8545 -5240
rect 5804 -5308 5900 -5292
rect 8816 -5292 8832 -2868
rect 8896 -5292 8912 -2868
rect 8816 -5308 8912 -5292
rect -6244 -5588 -6148 -5572
rect -8837 -5640 -6515 -5639
rect -8837 -7960 -8836 -5640
rect -6516 -7960 -6515 -5640
rect -8837 -7961 -6515 -7960
rect -6244 -8012 -6228 -5588
rect -6164 -8012 -6148 -5588
rect -3232 -5588 -3136 -5572
rect -5825 -5640 -3503 -5639
rect -5825 -7960 -5824 -5640
rect -3504 -7960 -3503 -5640
rect -5825 -7961 -3503 -7960
rect -6244 -8028 -6148 -8012
rect -3232 -8012 -3216 -5588
rect -3152 -8012 -3136 -5588
rect -220 -5588 -124 -5572
rect -2813 -5640 -491 -5639
rect -2813 -7960 -2812 -5640
rect -492 -7960 -491 -5640
rect -2813 -7961 -491 -7960
rect -3232 -8028 -3136 -8012
rect -220 -8012 -204 -5588
rect -140 -8012 -124 -5588
rect 2792 -5588 2888 -5572
rect 199 -5640 2521 -5639
rect 199 -7960 200 -5640
rect 2520 -7960 2521 -5640
rect 199 -7961 2521 -7960
rect -220 -8028 -124 -8012
rect 2792 -8012 2808 -5588
rect 2872 -8012 2888 -5588
rect 5804 -5588 5900 -5572
rect 3211 -5640 5533 -5639
rect 3211 -7960 3212 -5640
rect 5532 -7960 5533 -5640
rect 3211 -7961 5533 -7960
rect 2792 -8028 2888 -8012
rect 5804 -8012 5820 -5588
rect 5884 -8012 5900 -5588
rect 8816 -5588 8912 -5572
rect 6223 -5640 8545 -5639
rect 6223 -7960 6224 -5640
rect 8544 -7960 8545 -5640
rect 6223 -7961 8545 -7960
rect 5804 -8028 5900 -8012
rect 8816 -8012 8832 -5588
rect 8896 -8012 8912 -5588
rect 8816 -8028 8912 -8012
<< properties >>
string FIXED_BBOX 6144 5560 8624 8040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 12 l 12 val 297.12 carea 2.00 cperi 0.19 nx 6 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>

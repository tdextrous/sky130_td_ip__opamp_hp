magic
tech sky130A
magscale 1 2
timestamp 1714584774
<< error_p >>
rect -427 272 -363 278
rect -269 272 -205 278
rect -111 272 -47 278
rect 47 272 111 278
rect 205 272 269 278
rect 363 272 427 278
rect -427 238 -415 272
rect -269 238 -257 272
rect -111 238 -99 272
rect 47 238 59 272
rect 205 238 217 272
rect 363 238 375 272
rect -427 232 -363 238
rect -269 232 -205 238
rect -111 232 -47 238
rect 47 232 111 238
rect 205 232 269 238
rect 363 232 427 238
rect -427 -238 -363 -232
rect -269 -238 -205 -232
rect -111 -238 -47 -232
rect 47 -238 111 -232
rect 205 -238 269 -232
rect 363 -238 427 -232
rect -427 -272 -415 -238
rect -269 -272 -257 -238
rect -111 -272 -99 -238
rect 47 -272 59 -238
rect 205 -272 217 -238
rect 363 -272 375 -238
rect -427 -278 -363 -272
rect -269 -278 -205 -272
rect -111 -278 -47 -272
rect 47 -278 111 -272
rect 205 -278 269 -272
rect 363 -278 427 -272
<< pwell >>
rect -673 -458 673 458
<< mvnmos >>
rect -445 -200 -345 200
rect -287 -200 -187 200
rect -129 -200 -29 200
rect 29 -200 129 200
rect 187 -200 287 200
rect 345 -200 445 200
<< mvndiff >>
rect -503 188 -445 200
rect -503 -188 -491 188
rect -457 -188 -445 188
rect -503 -200 -445 -188
rect -345 188 -287 200
rect -345 -188 -333 188
rect -299 -188 -287 188
rect -345 -200 -287 -188
rect -187 188 -129 200
rect -187 -188 -175 188
rect -141 -188 -129 188
rect -187 -200 -129 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 129 188 187 200
rect 129 -188 141 188
rect 175 -188 187 188
rect 129 -200 187 -188
rect 287 188 345 200
rect 287 -188 299 188
rect 333 -188 345 188
rect 287 -200 345 -188
rect 445 188 503 200
rect 445 -188 457 188
rect 491 -188 503 188
rect 445 -200 503 -188
<< mvndiffc >>
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
<< mvpsubdiff >>
rect -637 410 637 422
rect -637 376 -529 410
rect 529 376 637 410
rect -637 364 637 376
rect -637 -364 -579 364
rect 579 -364 637 364
rect -637 -376 637 -364
rect -637 -410 -529 -376
rect 529 -410 637 -376
rect -637 -422 637 -410
<< mvpsubdiffcont >>
rect -529 376 529 410
rect -529 -410 529 -376
<< poly >>
rect -431 272 -359 288
rect -431 255 -415 272
rect -445 238 -415 255
rect -375 255 -359 272
rect -273 272 -201 288
rect -273 255 -257 272
rect -375 238 -345 255
rect -445 200 -345 238
rect -287 238 -257 255
rect -217 255 -201 272
rect -115 272 -43 288
rect -115 255 -99 272
rect -217 238 -187 255
rect -287 200 -187 238
rect -129 238 -99 255
rect -59 255 -43 272
rect 43 272 115 288
rect 43 255 59 272
rect -59 238 -29 255
rect -129 200 -29 238
rect 29 238 59 255
rect 99 255 115 272
rect 201 272 273 288
rect 201 255 217 272
rect 99 238 129 255
rect 29 200 129 238
rect 187 238 217 255
rect 257 255 273 272
rect 359 272 431 288
rect 359 255 375 272
rect 257 238 287 255
rect 187 200 287 238
rect 345 238 375 255
rect 415 255 431 272
rect 415 238 445 255
rect 345 200 445 238
rect -445 -238 -345 -200
rect -445 -255 -415 -238
rect -431 -272 -415 -255
rect -375 -255 -345 -238
rect -287 -238 -187 -200
rect -287 -255 -257 -238
rect -375 -272 -359 -255
rect -431 -288 -359 -272
rect -273 -272 -257 -255
rect -217 -255 -187 -238
rect -129 -238 -29 -200
rect -129 -255 -99 -238
rect -217 -272 -201 -255
rect -273 -288 -201 -272
rect -115 -272 -99 -255
rect -59 -255 -29 -238
rect 29 -238 129 -200
rect 29 -255 59 -238
rect -59 -272 -43 -255
rect -115 -288 -43 -272
rect 43 -272 59 -255
rect 99 -255 129 -238
rect 187 -238 287 -200
rect 187 -255 217 -238
rect 99 -272 115 -255
rect 43 -288 115 -272
rect 201 -272 217 -255
rect 257 -255 287 -238
rect 345 -238 445 -200
rect 345 -255 375 -238
rect 257 -272 273 -255
rect 201 -288 273 -272
rect 359 -272 375 -255
rect 415 -255 445 -238
rect 415 -272 431 -255
rect 359 -288 431 -272
<< polycont >>
rect -415 238 -375 272
rect -257 238 -217 272
rect -99 238 -59 272
rect 59 238 99 272
rect 217 238 257 272
rect 375 238 415 272
rect -415 -272 -375 -238
rect -257 -272 -217 -238
rect -99 -272 -59 -238
rect 59 -272 99 -238
rect 217 -272 257 -238
rect 375 -272 415 -238
<< locali >>
rect -625 376 -529 410
rect 529 376 625 410
rect -625 -376 -591 376
rect -431 238 -415 272
rect -375 238 -359 272
rect -273 238 -257 272
rect -217 238 -201 272
rect -115 238 -99 272
rect -59 238 -43 272
rect 43 238 59 272
rect 99 238 115 272
rect 201 238 217 272
rect 257 238 273 272
rect 359 238 375 272
rect 415 238 431 272
rect -491 188 -457 204
rect -491 -204 -457 -188
rect -333 188 -299 204
rect -333 -204 -299 -188
rect -175 188 -141 204
rect -175 -204 -141 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 141 188 175 204
rect 141 -204 175 -188
rect 299 188 333 204
rect 299 -204 333 -188
rect 457 188 491 204
rect 457 -204 491 -188
rect -431 -272 -415 -238
rect -375 -272 -359 -238
rect -273 -272 -257 -238
rect -217 -272 -201 -238
rect -115 -272 -99 -238
rect -59 -272 -43 -238
rect 43 -272 59 -238
rect 99 -272 115 -238
rect 201 -272 217 -238
rect 257 -272 273 -238
rect 359 -272 375 -238
rect 415 -272 431 -238
rect 591 -376 625 376
rect -625 -410 -529 -376
rect 529 -410 625 -376
<< viali >>
rect -415 238 -375 272
rect -257 238 -217 272
rect -99 238 -59 272
rect 59 238 99 272
rect 217 238 257 272
rect 375 238 415 272
rect -491 -188 -457 188
rect -333 -188 -299 188
rect -175 -188 -141 188
rect -17 -188 17 188
rect 141 -188 175 188
rect 299 -188 333 188
rect 457 -188 491 188
rect -415 -272 -375 -238
rect -257 -272 -217 -238
rect -99 -272 -59 -238
rect 59 -272 99 -238
rect 217 -272 257 -238
rect 375 -272 415 -238
<< metal1 >>
rect -427 272 -363 278
rect -427 238 -415 272
rect -375 238 -363 272
rect -427 232 -363 238
rect -269 272 -205 278
rect -269 238 -257 272
rect -217 238 -205 272
rect -269 232 -205 238
rect -111 272 -47 278
rect -111 238 -99 272
rect -59 238 -47 272
rect -111 232 -47 238
rect 47 272 111 278
rect 47 238 59 272
rect 99 238 111 272
rect 47 232 111 238
rect 205 272 269 278
rect 205 238 217 272
rect 257 238 269 272
rect 205 232 269 238
rect 363 272 427 278
rect 363 238 375 272
rect 415 238 427 272
rect 363 232 427 238
rect -497 188 -451 200
rect -497 -188 -491 188
rect -457 -188 -451 188
rect -497 -200 -451 -188
rect -339 188 -293 200
rect -339 -188 -333 188
rect -299 -188 -293 188
rect -339 -200 -293 -188
rect -181 188 -135 200
rect -181 -188 -175 188
rect -141 -188 -135 188
rect -181 -200 -135 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 135 188 181 200
rect 135 -188 141 188
rect 175 -188 181 188
rect 135 -200 181 -188
rect 293 188 339 200
rect 293 -188 299 188
rect 333 -188 339 188
rect 293 -200 339 -188
rect 451 188 497 200
rect 451 -188 457 188
rect 491 -188 497 188
rect 451 -200 497 -188
rect -427 -238 -363 -232
rect -427 -272 -415 -238
rect -375 -272 -363 -238
rect -427 -278 -363 -272
rect -269 -238 -205 -232
rect -269 -272 -257 -238
rect -217 -272 -205 -238
rect -269 -278 -205 -272
rect -111 -238 -47 -232
rect -111 -272 -99 -238
rect -59 -272 -47 -238
rect -111 -278 -47 -272
rect 47 -238 111 -232
rect 47 -272 59 -238
rect 99 -272 111 -238
rect 47 -278 111 -272
rect 205 -238 269 -232
rect 205 -272 217 -238
rect 257 -272 269 -238
rect 205 -278 269 -272
rect 363 -238 427 -232
rect 363 -272 375 -238
rect 415 -272 427 -238
rect 363 -278 427 -272
<< properties >>
string FIXED_BBOX -608 -393 608 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 6 diffcov 100 polycov 60 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713300419
<< pwell >>
rect -1876 -458 1876 458
<< mvnmos >>
rect -1648 -200 -1448 200
rect -1390 -200 -1190 200
rect -1132 -200 -932 200
rect -874 -200 -674 200
rect -616 -200 -416 200
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
rect 416 -200 616 200
rect 674 -200 874 200
rect 932 -200 1132 200
rect 1190 -200 1390 200
rect 1448 -200 1648 200
<< mvndiff >>
rect -1706 188 -1648 200
rect -1706 -188 -1694 188
rect -1660 -188 -1648 188
rect -1706 -200 -1648 -188
rect -1448 188 -1390 200
rect -1448 -188 -1436 188
rect -1402 -188 -1390 188
rect -1448 -200 -1390 -188
rect -1190 188 -1132 200
rect -1190 -188 -1178 188
rect -1144 -188 -1132 188
rect -1190 -200 -1132 -188
rect -932 188 -874 200
rect -932 -188 -920 188
rect -886 -188 -874 188
rect -932 -200 -874 -188
rect -674 188 -616 200
rect -674 -188 -662 188
rect -628 -188 -616 188
rect -674 -200 -616 -188
rect -416 188 -358 200
rect -416 -188 -404 188
rect -370 -188 -358 188
rect -416 -200 -358 -188
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
rect 358 188 416 200
rect 358 -188 370 188
rect 404 -188 416 188
rect 358 -200 416 -188
rect 616 188 674 200
rect 616 -188 628 188
rect 662 -188 674 188
rect 616 -200 674 -188
rect 874 188 932 200
rect 874 -188 886 188
rect 920 -188 932 188
rect 874 -200 932 -188
rect 1132 188 1190 200
rect 1132 -188 1144 188
rect 1178 -188 1190 188
rect 1132 -200 1190 -188
rect 1390 188 1448 200
rect 1390 -188 1402 188
rect 1436 -188 1448 188
rect 1390 -200 1448 -188
rect 1648 188 1706 200
rect 1648 -188 1660 188
rect 1694 -188 1706 188
rect 1648 -200 1706 -188
<< mvndiffc >>
rect -1694 -188 -1660 188
rect -1436 -188 -1402 188
rect -1178 -188 -1144 188
rect -920 -188 -886 188
rect -662 -188 -628 188
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect 628 -188 662 188
rect 886 -188 920 188
rect 1144 -188 1178 188
rect 1402 -188 1436 188
rect 1660 -188 1694 188
<< mvpsubdiff >>
rect -1840 410 1840 422
rect -1840 376 -1732 410
rect 1732 376 1840 410
rect -1840 364 1840 376
rect -1840 314 -1782 364
rect -1840 -314 -1828 314
rect -1794 -314 -1782 314
rect 1782 314 1840 364
rect -1840 -364 -1782 -314
rect 1782 -314 1794 314
rect 1828 -314 1840 314
rect 1782 -364 1840 -314
rect -1840 -376 1840 -364
rect -1840 -410 -1732 -376
rect 1732 -410 1840 -376
rect -1840 -422 1840 -410
<< mvpsubdiffcont >>
rect -1732 376 1732 410
rect -1828 -314 -1794 314
rect 1794 -314 1828 314
rect -1732 -410 1732 -376
<< poly >>
rect -1614 272 -1482 288
rect -1614 255 -1598 272
rect -1648 238 -1598 255
rect -1498 255 -1482 272
rect -1356 272 -1224 288
rect -1356 255 -1340 272
rect -1498 238 -1448 255
rect -1648 200 -1448 238
rect -1390 238 -1340 255
rect -1240 255 -1224 272
rect -1098 272 -966 288
rect -1098 255 -1082 272
rect -1240 238 -1190 255
rect -1390 200 -1190 238
rect -1132 238 -1082 255
rect -982 255 -966 272
rect -840 272 -708 288
rect -840 255 -824 272
rect -982 238 -932 255
rect -1132 200 -932 238
rect -874 238 -824 255
rect -724 255 -708 272
rect -582 272 -450 288
rect -582 255 -566 272
rect -724 238 -674 255
rect -874 200 -674 238
rect -616 238 -566 255
rect -466 255 -450 272
rect -324 272 -192 288
rect -324 255 -308 272
rect -466 238 -416 255
rect -616 200 -416 238
rect -358 238 -308 255
rect -208 255 -192 272
rect -66 272 66 288
rect -66 255 -50 272
rect -208 238 -158 255
rect -358 200 -158 238
rect -100 238 -50 255
rect 50 255 66 272
rect 192 272 324 288
rect 192 255 208 272
rect 50 238 100 255
rect -100 200 100 238
rect 158 238 208 255
rect 308 255 324 272
rect 450 272 582 288
rect 450 255 466 272
rect 308 238 358 255
rect 158 200 358 238
rect 416 238 466 255
rect 566 255 582 272
rect 708 272 840 288
rect 708 255 724 272
rect 566 238 616 255
rect 416 200 616 238
rect 674 238 724 255
rect 824 255 840 272
rect 966 272 1098 288
rect 966 255 982 272
rect 824 238 874 255
rect 674 200 874 238
rect 932 238 982 255
rect 1082 255 1098 272
rect 1224 272 1356 288
rect 1224 255 1240 272
rect 1082 238 1132 255
rect 932 200 1132 238
rect 1190 238 1240 255
rect 1340 255 1356 272
rect 1482 272 1614 288
rect 1482 255 1498 272
rect 1340 238 1390 255
rect 1190 200 1390 238
rect 1448 238 1498 255
rect 1598 255 1614 272
rect 1598 238 1648 255
rect 1448 200 1648 238
rect -1648 -238 -1448 -200
rect -1648 -255 -1598 -238
rect -1614 -272 -1598 -255
rect -1498 -255 -1448 -238
rect -1390 -238 -1190 -200
rect -1390 -255 -1340 -238
rect -1498 -272 -1482 -255
rect -1614 -288 -1482 -272
rect -1356 -272 -1340 -255
rect -1240 -255 -1190 -238
rect -1132 -238 -932 -200
rect -1132 -255 -1082 -238
rect -1240 -272 -1224 -255
rect -1356 -288 -1224 -272
rect -1098 -272 -1082 -255
rect -982 -255 -932 -238
rect -874 -238 -674 -200
rect -874 -255 -824 -238
rect -982 -272 -966 -255
rect -1098 -288 -966 -272
rect -840 -272 -824 -255
rect -724 -255 -674 -238
rect -616 -238 -416 -200
rect -616 -255 -566 -238
rect -724 -272 -708 -255
rect -840 -288 -708 -272
rect -582 -272 -566 -255
rect -466 -255 -416 -238
rect -358 -238 -158 -200
rect -358 -255 -308 -238
rect -466 -272 -450 -255
rect -582 -288 -450 -272
rect -324 -272 -308 -255
rect -208 -255 -158 -238
rect -100 -238 100 -200
rect -100 -255 -50 -238
rect -208 -272 -192 -255
rect -324 -288 -192 -272
rect -66 -272 -50 -255
rect 50 -255 100 -238
rect 158 -238 358 -200
rect 158 -255 208 -238
rect 50 -272 66 -255
rect -66 -288 66 -272
rect 192 -272 208 -255
rect 308 -255 358 -238
rect 416 -238 616 -200
rect 416 -255 466 -238
rect 308 -272 324 -255
rect 192 -288 324 -272
rect 450 -272 466 -255
rect 566 -255 616 -238
rect 674 -238 874 -200
rect 674 -255 724 -238
rect 566 -272 582 -255
rect 450 -288 582 -272
rect 708 -272 724 -255
rect 824 -255 874 -238
rect 932 -238 1132 -200
rect 932 -255 982 -238
rect 824 -272 840 -255
rect 708 -288 840 -272
rect 966 -272 982 -255
rect 1082 -255 1132 -238
rect 1190 -238 1390 -200
rect 1190 -255 1240 -238
rect 1082 -272 1098 -255
rect 966 -288 1098 -272
rect 1224 -272 1240 -255
rect 1340 -255 1390 -238
rect 1448 -238 1648 -200
rect 1448 -255 1498 -238
rect 1340 -272 1356 -255
rect 1224 -288 1356 -272
rect 1482 -272 1498 -255
rect 1598 -255 1648 -238
rect 1598 -272 1614 -255
rect 1482 -288 1614 -272
<< polycont >>
rect -1598 238 -1498 272
rect -1340 238 -1240 272
rect -1082 238 -982 272
rect -824 238 -724 272
rect -566 238 -466 272
rect -308 238 -208 272
rect -50 238 50 272
rect 208 238 308 272
rect 466 238 566 272
rect 724 238 824 272
rect 982 238 1082 272
rect 1240 238 1340 272
rect 1498 238 1598 272
rect -1598 -272 -1498 -238
rect -1340 -272 -1240 -238
rect -1082 -272 -982 -238
rect -824 -272 -724 -238
rect -566 -272 -466 -238
rect -308 -272 -208 -238
rect -50 -272 50 -238
rect 208 -272 308 -238
rect 466 -272 566 -238
rect 724 -272 824 -238
rect 982 -272 1082 -238
rect 1240 -272 1340 -238
rect 1498 -272 1598 -238
<< locali >>
rect -1828 376 -1732 410
rect 1732 376 1828 410
rect -1828 314 -1794 376
rect 1794 314 1828 376
rect -1614 238 -1598 272
rect -1498 238 -1482 272
rect -1356 238 -1340 272
rect -1240 238 -1224 272
rect -1098 238 -1082 272
rect -982 238 -966 272
rect -840 238 -824 272
rect -724 238 -708 272
rect -582 238 -566 272
rect -466 238 -450 272
rect -324 238 -308 272
rect -208 238 -192 272
rect -66 238 -50 272
rect 50 238 66 272
rect 192 238 208 272
rect 308 238 324 272
rect 450 238 466 272
rect 566 238 582 272
rect 708 238 724 272
rect 824 238 840 272
rect 966 238 982 272
rect 1082 238 1098 272
rect 1224 238 1240 272
rect 1340 238 1356 272
rect 1482 238 1498 272
rect 1598 238 1614 272
rect -1694 188 -1660 204
rect -1694 -204 -1660 -188
rect -1436 188 -1402 204
rect -1436 -204 -1402 -188
rect -1178 188 -1144 204
rect -1178 -204 -1144 -188
rect -920 188 -886 204
rect -920 -204 -886 -188
rect -662 188 -628 204
rect -662 -204 -628 -188
rect -404 188 -370 204
rect -404 -204 -370 -188
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect 370 188 404 204
rect 370 -204 404 -188
rect 628 188 662 204
rect 628 -204 662 -188
rect 886 188 920 204
rect 886 -204 920 -188
rect 1144 188 1178 204
rect 1144 -204 1178 -188
rect 1402 188 1436 204
rect 1402 -204 1436 -188
rect 1660 188 1694 204
rect 1660 -204 1694 -188
rect -1614 -272 -1598 -238
rect -1498 -272 -1482 -238
rect -1356 -272 -1340 -238
rect -1240 -272 -1224 -238
rect -1098 -272 -1082 -238
rect -982 -272 -966 -238
rect -840 -272 -824 -238
rect -724 -272 -708 -238
rect -582 -272 -566 -238
rect -466 -272 -450 -238
rect -324 -272 -308 -238
rect -208 -272 -192 -238
rect -66 -272 -50 -238
rect 50 -272 66 -238
rect 192 -272 208 -238
rect 308 -272 324 -238
rect 450 -272 466 -238
rect 566 -272 582 -238
rect 708 -272 724 -238
rect 824 -272 840 -238
rect 966 -272 982 -238
rect 1082 -272 1098 -238
rect 1224 -272 1240 -238
rect 1340 -272 1356 -238
rect 1482 -272 1498 -238
rect 1598 -272 1614 -238
rect -1828 -376 -1794 -314
rect 1794 -376 1828 -314
rect -1828 -410 -1732 -376
rect 1732 -410 1828 -376
<< viali >>
rect -1598 238 -1498 272
rect -1340 238 -1240 272
rect -1082 238 -982 272
rect -824 238 -724 272
rect -566 238 -466 272
rect -308 238 -208 272
rect -50 238 50 272
rect 208 238 308 272
rect 466 238 566 272
rect 724 238 824 272
rect 982 238 1082 272
rect 1240 238 1340 272
rect 1498 238 1598 272
rect -1694 -188 -1660 188
rect -1436 -188 -1402 188
rect -1178 -188 -1144 188
rect -920 -188 -886 188
rect -662 -188 -628 188
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect 628 -188 662 188
rect 886 -188 920 188
rect 1144 -188 1178 188
rect 1402 -188 1436 188
rect 1660 -188 1694 188
rect -1598 -272 -1498 -238
rect -1340 -272 -1240 -238
rect -1082 -272 -982 -238
rect -824 -272 -724 -238
rect -566 -272 -466 -238
rect -308 -272 -208 -238
rect -50 -272 50 -238
rect 208 -272 308 -238
rect 466 -272 566 -238
rect 724 -272 824 -238
rect 982 -272 1082 -238
rect 1240 -272 1340 -238
rect 1498 -272 1598 -238
<< metal1 >>
rect -1610 272 -1486 278
rect -1610 238 -1598 272
rect -1498 238 -1486 272
rect -1610 232 -1486 238
rect -1352 272 -1228 278
rect -1352 238 -1340 272
rect -1240 238 -1228 272
rect -1352 232 -1228 238
rect -1094 272 -970 278
rect -1094 238 -1082 272
rect -982 238 -970 272
rect -1094 232 -970 238
rect -836 272 -712 278
rect -836 238 -824 272
rect -724 238 -712 272
rect -836 232 -712 238
rect -578 272 -454 278
rect -578 238 -566 272
rect -466 238 -454 272
rect -578 232 -454 238
rect -320 272 -196 278
rect -320 238 -308 272
rect -208 238 -196 272
rect -320 232 -196 238
rect -62 272 62 278
rect -62 238 -50 272
rect 50 238 62 272
rect -62 232 62 238
rect 196 272 320 278
rect 196 238 208 272
rect 308 238 320 272
rect 196 232 320 238
rect 454 272 578 278
rect 454 238 466 272
rect 566 238 578 272
rect 454 232 578 238
rect 712 272 836 278
rect 712 238 724 272
rect 824 238 836 272
rect 712 232 836 238
rect 970 272 1094 278
rect 970 238 982 272
rect 1082 238 1094 272
rect 970 232 1094 238
rect 1228 272 1352 278
rect 1228 238 1240 272
rect 1340 238 1352 272
rect 1228 232 1352 238
rect 1486 272 1610 278
rect 1486 238 1498 272
rect 1598 238 1610 272
rect 1486 232 1610 238
rect -1700 188 -1654 200
rect -1700 -188 -1694 188
rect -1660 -188 -1654 188
rect -1700 -200 -1654 -188
rect -1442 188 -1396 200
rect -1442 -188 -1436 188
rect -1402 -188 -1396 188
rect -1442 -200 -1396 -188
rect -1184 188 -1138 200
rect -1184 -188 -1178 188
rect -1144 -188 -1138 188
rect -1184 -200 -1138 -188
rect -926 188 -880 200
rect -926 -188 -920 188
rect -886 -188 -880 188
rect -926 -200 -880 -188
rect -668 188 -622 200
rect -668 -188 -662 188
rect -628 -188 -622 188
rect -668 -200 -622 -188
rect -410 188 -364 200
rect -410 -188 -404 188
rect -370 -188 -364 188
rect -410 -200 -364 -188
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect 364 188 410 200
rect 364 -188 370 188
rect 404 -188 410 188
rect 364 -200 410 -188
rect 622 188 668 200
rect 622 -188 628 188
rect 662 -188 668 188
rect 622 -200 668 -188
rect 880 188 926 200
rect 880 -188 886 188
rect 920 -188 926 188
rect 880 -200 926 -188
rect 1138 188 1184 200
rect 1138 -188 1144 188
rect 1178 -188 1184 188
rect 1138 -200 1184 -188
rect 1396 188 1442 200
rect 1396 -188 1402 188
rect 1436 -188 1442 188
rect 1396 -200 1442 -188
rect 1654 188 1700 200
rect 1654 -188 1660 188
rect 1694 -188 1700 188
rect 1654 -200 1700 -188
rect -1610 -238 -1486 -232
rect -1610 -272 -1598 -238
rect -1498 -272 -1486 -238
rect -1610 -278 -1486 -272
rect -1352 -238 -1228 -232
rect -1352 -272 -1340 -238
rect -1240 -272 -1228 -238
rect -1352 -278 -1228 -272
rect -1094 -238 -970 -232
rect -1094 -272 -1082 -238
rect -982 -272 -970 -238
rect -1094 -278 -970 -272
rect -836 -238 -712 -232
rect -836 -272 -824 -238
rect -724 -272 -712 -238
rect -836 -278 -712 -272
rect -578 -238 -454 -232
rect -578 -272 -566 -238
rect -466 -272 -454 -238
rect -578 -278 -454 -272
rect -320 -238 -196 -232
rect -320 -272 -308 -238
rect -208 -272 -196 -238
rect -320 -278 -196 -272
rect -62 -238 62 -232
rect -62 -272 -50 -238
rect 50 -272 62 -238
rect -62 -278 62 -272
rect 196 -238 320 -232
rect 196 -272 208 -238
rect 308 -272 320 -238
rect 196 -278 320 -272
rect 454 -238 578 -232
rect 454 -272 466 -238
rect 566 -272 578 -238
rect 454 -278 578 -272
rect 712 -238 836 -232
rect 712 -272 724 -238
rect 824 -272 836 -238
rect 712 -278 836 -272
rect 970 -238 1094 -232
rect 970 -272 982 -238
rect 1082 -272 1094 -238
rect 970 -278 1094 -272
rect 1228 -238 1352 -232
rect 1228 -272 1240 -238
rect 1340 -272 1352 -238
rect 1228 -278 1352 -272
rect 1486 -238 1610 -232
rect 1486 -272 1498 -238
rect 1598 -272 1610 -238
rect 1486 -278 1610 -272
<< properties >>
string FIXED_BBOX -1811 -393 1811 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 13 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

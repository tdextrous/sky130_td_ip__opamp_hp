magic
tech sky130A
magscale 1 2
timestamp 1713235147
<< pwell >>
rect -633 -1096 633 1096
<< psubdiff >>
rect -597 1026 -501 1060
rect 501 1026 597 1060
rect -597 964 -563 1026
rect 563 964 597 1026
rect -597 -1026 -563 -964
rect 563 -1026 597 -964
rect -597 -1060 -501 -1026
rect 501 -1060 597 -1026
<< psubdiffcont >>
rect -501 1026 501 1060
rect -597 -964 -563 964
rect 563 -964 597 964
rect -501 -1060 501 -1026
<< poly >>
rect -467 914 -387 930
rect -467 880 -451 914
rect -403 880 -387 914
rect -467 500 -387 880
rect -467 -880 -387 -500
rect -467 -914 -451 -880
rect -403 -914 -387 -880
rect -467 -930 -387 -914
rect -345 914 -265 930
rect -345 880 -329 914
rect -281 880 -265 914
rect -345 500 -265 880
rect -345 -880 -265 -500
rect -345 -914 -329 -880
rect -281 -914 -265 -880
rect -345 -930 -265 -914
rect -223 914 -143 930
rect -223 880 -207 914
rect -159 880 -143 914
rect -223 500 -143 880
rect -223 -880 -143 -500
rect -223 -914 -207 -880
rect -159 -914 -143 -880
rect -223 -930 -143 -914
rect -101 914 -21 930
rect -101 880 -85 914
rect -37 880 -21 914
rect -101 500 -21 880
rect -101 -880 -21 -500
rect -101 -914 -85 -880
rect -37 -914 -21 -880
rect -101 -930 -21 -914
rect 21 914 101 930
rect 21 880 37 914
rect 85 880 101 914
rect 21 500 101 880
rect 21 -880 101 -500
rect 21 -914 37 -880
rect 85 -914 101 -880
rect 21 -930 101 -914
rect 143 914 223 930
rect 143 880 159 914
rect 207 880 223 914
rect 143 500 223 880
rect 143 -880 223 -500
rect 143 -914 159 -880
rect 207 -914 223 -880
rect 143 -930 223 -914
rect 265 914 345 930
rect 265 880 281 914
rect 329 880 345 914
rect 265 500 345 880
rect 265 -880 345 -500
rect 265 -914 281 -880
rect 329 -914 345 -880
rect 265 -930 345 -914
rect 387 914 467 930
rect 387 880 403 914
rect 451 880 467 914
rect 387 500 467 880
rect 387 -880 467 -500
rect 387 -914 403 -880
rect 451 -914 467 -880
rect 387 -930 467 -914
<< polycont >>
rect -451 880 -403 914
rect -451 -914 -403 -880
rect -329 880 -281 914
rect -329 -914 -281 -880
rect -207 880 -159 914
rect -207 -914 -159 -880
rect -85 880 -37 914
rect -85 -914 -37 -880
rect 37 880 85 914
rect 37 -914 85 -880
rect 159 880 207 914
rect 159 -914 207 -880
rect 281 880 329 914
rect 281 -914 329 -880
rect 403 880 451 914
rect 403 -914 451 -880
<< npolyres >>
rect -467 -500 -387 500
rect -345 -500 -265 500
rect -223 -500 -143 500
rect -101 -500 -21 500
rect 21 -500 101 500
rect 143 -500 223 500
rect 265 -500 345 500
rect 387 -500 467 500
<< locali >>
rect -597 1026 -501 1060
rect 501 1026 597 1060
rect -597 964 -563 1026
rect 563 964 597 1026
rect -467 880 -451 914
rect -403 880 -387 914
rect -345 880 -329 914
rect -281 880 -265 914
rect -223 880 -207 914
rect -159 880 -143 914
rect -101 880 -85 914
rect -37 880 -21 914
rect 21 880 37 914
rect 85 880 101 914
rect 143 880 159 914
rect 207 880 223 914
rect 265 880 281 914
rect 329 880 345 914
rect 387 880 403 914
rect 451 880 467 914
rect -467 -914 -451 -880
rect -403 -914 -387 -880
rect -345 -914 -329 -880
rect -281 -914 -265 -880
rect -223 -914 -207 -880
rect -159 -914 -143 -880
rect -101 -914 -85 -880
rect -37 -914 -21 -880
rect 21 -914 37 -880
rect 85 -914 101 -880
rect 143 -914 159 -880
rect 207 -914 223 -880
rect 265 -914 281 -880
rect 329 -914 345 -880
rect 387 -914 403 -880
rect 451 -914 467 -880
rect -597 -1026 -563 -964
rect 563 -1026 597 -964
rect -597 -1060 -501 -1026
rect 501 -1060 597 -1026
<< viali >>
rect -451 880 -403 914
rect -329 880 -281 914
rect -207 880 -159 914
rect -85 880 -37 914
rect 37 880 85 914
rect 159 880 207 914
rect 281 880 329 914
rect 403 880 451 914
rect -451 517 -403 880
rect -329 517 -281 880
rect -207 517 -159 880
rect -85 517 -37 880
rect 37 517 85 880
rect 159 517 207 880
rect 281 517 329 880
rect 403 517 451 880
rect -451 -880 -403 -517
rect -329 -880 -281 -517
rect -207 -880 -159 -517
rect -85 -880 -37 -517
rect 37 -880 85 -517
rect 159 -880 207 -517
rect 281 -880 329 -517
rect 403 -880 451 -517
rect -451 -914 -403 -880
rect -329 -914 -281 -880
rect -207 -914 -159 -880
rect -85 -914 -37 -880
rect 37 -914 85 -880
rect 159 -914 207 -880
rect 281 -914 329 -880
rect 403 -914 451 -880
<< metal1 >>
rect -457 914 -397 926
rect -457 517 -451 914
rect -403 517 -397 914
rect -457 505 -397 517
rect -335 914 -275 926
rect -335 517 -329 914
rect -281 517 -275 914
rect -335 505 -275 517
rect -213 914 -153 926
rect -213 517 -207 914
rect -159 517 -153 914
rect -213 505 -153 517
rect -91 914 -31 926
rect -91 517 -85 914
rect -37 517 -31 914
rect -91 505 -31 517
rect 31 914 91 926
rect 31 517 37 914
rect 85 517 91 914
rect 31 505 91 517
rect 153 914 213 926
rect 153 517 159 914
rect 207 517 213 914
rect 153 505 213 517
rect 275 914 335 926
rect 275 517 281 914
rect 329 517 335 914
rect 275 505 335 517
rect 397 914 457 926
rect 397 517 403 914
rect 451 517 457 914
rect 397 505 457 517
rect -457 -517 -397 -505
rect -457 -914 -451 -517
rect -403 -914 -397 -517
rect -457 -926 -397 -914
rect -335 -517 -275 -505
rect -335 -914 -329 -517
rect -281 -914 -275 -517
rect -335 -926 -275 -914
rect -213 -517 -153 -505
rect -213 -914 -207 -517
rect -159 -914 -153 -517
rect -213 -926 -153 -914
rect -91 -517 -31 -505
rect -91 -914 -85 -517
rect -37 -914 -31 -517
rect -91 -926 -31 -914
rect 31 -517 91 -505
rect 31 -914 37 -517
rect 85 -914 91 -517
rect 31 -926 91 -914
rect 153 -517 213 -505
rect 153 -914 159 -517
rect 207 -914 213 -517
rect 153 -926 213 -914
rect 275 -517 335 -505
rect 275 -914 281 -517
rect 329 -914 335 -517
rect 275 -926 335 -914
rect 397 -517 457 -505
rect 397 -914 403 -517
rect 451 -914 457 -517
rect 397 -926 457 -914
<< properties >>
string FIXED_BBOX -580 -1043 580 1043
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.4 l 5 m 1 nx 8 wmin 0.330 lmin 1.650 rho 48.2 val 602.5 dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

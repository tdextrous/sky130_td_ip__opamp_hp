magic
tech sky130A
magscale 1 2
timestamp 1713233716
<< nwell >>
rect -4357 -697 4357 697
<< mvpmos >>
rect -4099 -400 -3899 400
rect -3841 -400 -3641 400
rect -3583 -400 -3383 400
rect -3325 -400 -3125 400
rect -3067 -400 -2867 400
rect -2809 -400 -2609 400
rect -2551 -400 -2351 400
rect -2293 -400 -2093 400
rect -2035 -400 -1835 400
rect -1777 -400 -1577 400
rect -1519 -400 -1319 400
rect -1261 -400 -1061 400
rect -1003 -400 -803 400
rect -745 -400 -545 400
rect -487 -400 -287 400
rect -229 -400 -29 400
rect 29 -400 229 400
rect 287 -400 487 400
rect 545 -400 745 400
rect 803 -400 1003 400
rect 1061 -400 1261 400
rect 1319 -400 1519 400
rect 1577 -400 1777 400
rect 1835 -400 2035 400
rect 2093 -400 2293 400
rect 2351 -400 2551 400
rect 2609 -400 2809 400
rect 2867 -400 3067 400
rect 3125 -400 3325 400
rect 3383 -400 3583 400
rect 3641 -400 3841 400
rect 3899 -400 4099 400
<< mvpdiff >>
rect -4157 388 -4099 400
rect -4157 -388 -4145 388
rect -4111 -388 -4099 388
rect -4157 -400 -4099 -388
rect -3899 388 -3841 400
rect -3899 -388 -3887 388
rect -3853 -388 -3841 388
rect -3899 -400 -3841 -388
rect -3641 388 -3583 400
rect -3641 -388 -3629 388
rect -3595 -388 -3583 388
rect -3641 -400 -3583 -388
rect -3383 388 -3325 400
rect -3383 -388 -3371 388
rect -3337 -388 -3325 388
rect -3383 -400 -3325 -388
rect -3125 388 -3067 400
rect -3125 -388 -3113 388
rect -3079 -388 -3067 388
rect -3125 -400 -3067 -388
rect -2867 388 -2809 400
rect -2867 -388 -2855 388
rect -2821 -388 -2809 388
rect -2867 -400 -2809 -388
rect -2609 388 -2551 400
rect -2609 -388 -2597 388
rect -2563 -388 -2551 388
rect -2609 -400 -2551 -388
rect -2351 388 -2293 400
rect -2351 -388 -2339 388
rect -2305 -388 -2293 388
rect -2351 -400 -2293 -388
rect -2093 388 -2035 400
rect -2093 -388 -2081 388
rect -2047 -388 -2035 388
rect -2093 -400 -2035 -388
rect -1835 388 -1777 400
rect -1835 -388 -1823 388
rect -1789 -388 -1777 388
rect -1835 -400 -1777 -388
rect -1577 388 -1519 400
rect -1577 -388 -1565 388
rect -1531 -388 -1519 388
rect -1577 -400 -1519 -388
rect -1319 388 -1261 400
rect -1319 -388 -1307 388
rect -1273 -388 -1261 388
rect -1319 -400 -1261 -388
rect -1061 388 -1003 400
rect -1061 -388 -1049 388
rect -1015 -388 -1003 388
rect -1061 -400 -1003 -388
rect -803 388 -745 400
rect -803 -388 -791 388
rect -757 -388 -745 388
rect -803 -400 -745 -388
rect -545 388 -487 400
rect -545 -388 -533 388
rect -499 -388 -487 388
rect -545 -400 -487 -388
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
rect 487 388 545 400
rect 487 -388 499 388
rect 533 -388 545 388
rect 487 -400 545 -388
rect 745 388 803 400
rect 745 -388 757 388
rect 791 -388 803 388
rect 745 -400 803 -388
rect 1003 388 1061 400
rect 1003 -388 1015 388
rect 1049 -388 1061 388
rect 1003 -400 1061 -388
rect 1261 388 1319 400
rect 1261 -388 1273 388
rect 1307 -388 1319 388
rect 1261 -400 1319 -388
rect 1519 388 1577 400
rect 1519 -388 1531 388
rect 1565 -388 1577 388
rect 1519 -400 1577 -388
rect 1777 388 1835 400
rect 1777 -388 1789 388
rect 1823 -388 1835 388
rect 1777 -400 1835 -388
rect 2035 388 2093 400
rect 2035 -388 2047 388
rect 2081 -388 2093 388
rect 2035 -400 2093 -388
rect 2293 388 2351 400
rect 2293 -388 2305 388
rect 2339 -388 2351 388
rect 2293 -400 2351 -388
rect 2551 388 2609 400
rect 2551 -388 2563 388
rect 2597 -388 2609 388
rect 2551 -400 2609 -388
rect 2809 388 2867 400
rect 2809 -388 2821 388
rect 2855 -388 2867 388
rect 2809 -400 2867 -388
rect 3067 388 3125 400
rect 3067 -388 3079 388
rect 3113 -388 3125 388
rect 3067 -400 3125 -388
rect 3325 388 3383 400
rect 3325 -388 3337 388
rect 3371 -388 3383 388
rect 3325 -400 3383 -388
rect 3583 388 3641 400
rect 3583 -388 3595 388
rect 3629 -388 3641 388
rect 3583 -400 3641 -388
rect 3841 388 3899 400
rect 3841 -388 3853 388
rect 3887 -388 3899 388
rect 3841 -400 3899 -388
rect 4099 388 4157 400
rect 4099 -388 4111 388
rect 4145 -388 4157 388
rect 4099 -400 4157 -388
<< mvpdiffc >>
rect -4145 -388 -4111 388
rect -3887 -388 -3853 388
rect -3629 -388 -3595 388
rect -3371 -388 -3337 388
rect -3113 -388 -3079 388
rect -2855 -388 -2821 388
rect -2597 -388 -2563 388
rect -2339 -388 -2305 388
rect -2081 -388 -2047 388
rect -1823 -388 -1789 388
rect -1565 -388 -1531 388
rect -1307 -388 -1273 388
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect 1273 -388 1307 388
rect 1531 -388 1565 388
rect 1789 -388 1823 388
rect 2047 -388 2081 388
rect 2305 -388 2339 388
rect 2563 -388 2597 388
rect 2821 -388 2855 388
rect 3079 -388 3113 388
rect 3337 -388 3371 388
rect 3595 -388 3629 388
rect 3853 -388 3887 388
rect 4111 -388 4145 388
<< mvnsubdiff >>
rect -4291 619 4291 631
rect -4291 585 -4183 619
rect 4183 585 4291 619
rect -4291 573 4291 585
rect -4291 523 -4233 573
rect -4291 -523 -4279 523
rect -4245 -523 -4233 523
rect 4233 523 4291 573
rect -4291 -573 -4233 -523
rect 4233 -523 4245 523
rect 4279 -523 4291 523
rect 4233 -573 4291 -523
rect -4291 -585 4291 -573
rect -4291 -619 -4183 -585
rect 4183 -619 4291 -585
rect -4291 -631 4291 -619
<< mvnsubdiffcont >>
rect -4183 585 4183 619
rect -4279 -523 -4245 523
rect 4245 -523 4279 523
rect -4183 -619 4183 -585
<< poly >>
rect -4099 481 -3899 497
rect -4099 447 -4083 481
rect -3915 447 -3899 481
rect -4099 400 -3899 447
rect -3841 481 -3641 497
rect -3841 447 -3825 481
rect -3657 447 -3641 481
rect -3841 400 -3641 447
rect -3583 481 -3383 497
rect -3583 447 -3567 481
rect -3399 447 -3383 481
rect -3583 400 -3383 447
rect -3325 481 -3125 497
rect -3325 447 -3309 481
rect -3141 447 -3125 481
rect -3325 400 -3125 447
rect -3067 481 -2867 497
rect -3067 447 -3051 481
rect -2883 447 -2867 481
rect -3067 400 -2867 447
rect -2809 481 -2609 497
rect -2809 447 -2793 481
rect -2625 447 -2609 481
rect -2809 400 -2609 447
rect -2551 481 -2351 497
rect -2551 447 -2535 481
rect -2367 447 -2351 481
rect -2551 400 -2351 447
rect -2293 481 -2093 497
rect -2293 447 -2277 481
rect -2109 447 -2093 481
rect -2293 400 -2093 447
rect -2035 481 -1835 497
rect -2035 447 -2019 481
rect -1851 447 -1835 481
rect -2035 400 -1835 447
rect -1777 481 -1577 497
rect -1777 447 -1761 481
rect -1593 447 -1577 481
rect -1777 400 -1577 447
rect -1519 481 -1319 497
rect -1519 447 -1503 481
rect -1335 447 -1319 481
rect -1519 400 -1319 447
rect -1261 481 -1061 497
rect -1261 447 -1245 481
rect -1077 447 -1061 481
rect -1261 400 -1061 447
rect -1003 481 -803 497
rect -1003 447 -987 481
rect -819 447 -803 481
rect -1003 400 -803 447
rect -745 481 -545 497
rect -745 447 -729 481
rect -561 447 -545 481
rect -745 400 -545 447
rect -487 481 -287 497
rect -487 447 -471 481
rect -303 447 -287 481
rect -487 400 -287 447
rect -229 481 -29 497
rect -229 447 -213 481
rect -45 447 -29 481
rect -229 400 -29 447
rect 29 481 229 497
rect 29 447 45 481
rect 213 447 229 481
rect 29 400 229 447
rect 287 481 487 497
rect 287 447 303 481
rect 471 447 487 481
rect 287 400 487 447
rect 545 481 745 497
rect 545 447 561 481
rect 729 447 745 481
rect 545 400 745 447
rect 803 481 1003 497
rect 803 447 819 481
rect 987 447 1003 481
rect 803 400 1003 447
rect 1061 481 1261 497
rect 1061 447 1077 481
rect 1245 447 1261 481
rect 1061 400 1261 447
rect 1319 481 1519 497
rect 1319 447 1335 481
rect 1503 447 1519 481
rect 1319 400 1519 447
rect 1577 481 1777 497
rect 1577 447 1593 481
rect 1761 447 1777 481
rect 1577 400 1777 447
rect 1835 481 2035 497
rect 1835 447 1851 481
rect 2019 447 2035 481
rect 1835 400 2035 447
rect 2093 481 2293 497
rect 2093 447 2109 481
rect 2277 447 2293 481
rect 2093 400 2293 447
rect 2351 481 2551 497
rect 2351 447 2367 481
rect 2535 447 2551 481
rect 2351 400 2551 447
rect 2609 481 2809 497
rect 2609 447 2625 481
rect 2793 447 2809 481
rect 2609 400 2809 447
rect 2867 481 3067 497
rect 2867 447 2883 481
rect 3051 447 3067 481
rect 2867 400 3067 447
rect 3125 481 3325 497
rect 3125 447 3141 481
rect 3309 447 3325 481
rect 3125 400 3325 447
rect 3383 481 3583 497
rect 3383 447 3399 481
rect 3567 447 3583 481
rect 3383 400 3583 447
rect 3641 481 3841 497
rect 3641 447 3657 481
rect 3825 447 3841 481
rect 3641 400 3841 447
rect 3899 481 4099 497
rect 3899 447 3915 481
rect 4083 447 4099 481
rect 3899 400 4099 447
rect -4099 -447 -3899 -400
rect -4099 -481 -4083 -447
rect -3915 -481 -3899 -447
rect -4099 -497 -3899 -481
rect -3841 -447 -3641 -400
rect -3841 -481 -3825 -447
rect -3657 -481 -3641 -447
rect -3841 -497 -3641 -481
rect -3583 -447 -3383 -400
rect -3583 -481 -3567 -447
rect -3399 -481 -3383 -447
rect -3583 -497 -3383 -481
rect -3325 -447 -3125 -400
rect -3325 -481 -3309 -447
rect -3141 -481 -3125 -447
rect -3325 -497 -3125 -481
rect -3067 -447 -2867 -400
rect -3067 -481 -3051 -447
rect -2883 -481 -2867 -447
rect -3067 -497 -2867 -481
rect -2809 -447 -2609 -400
rect -2809 -481 -2793 -447
rect -2625 -481 -2609 -447
rect -2809 -497 -2609 -481
rect -2551 -447 -2351 -400
rect -2551 -481 -2535 -447
rect -2367 -481 -2351 -447
rect -2551 -497 -2351 -481
rect -2293 -447 -2093 -400
rect -2293 -481 -2277 -447
rect -2109 -481 -2093 -447
rect -2293 -497 -2093 -481
rect -2035 -447 -1835 -400
rect -2035 -481 -2019 -447
rect -1851 -481 -1835 -447
rect -2035 -497 -1835 -481
rect -1777 -447 -1577 -400
rect -1777 -481 -1761 -447
rect -1593 -481 -1577 -447
rect -1777 -497 -1577 -481
rect -1519 -447 -1319 -400
rect -1519 -481 -1503 -447
rect -1335 -481 -1319 -447
rect -1519 -497 -1319 -481
rect -1261 -447 -1061 -400
rect -1261 -481 -1245 -447
rect -1077 -481 -1061 -447
rect -1261 -497 -1061 -481
rect -1003 -447 -803 -400
rect -1003 -481 -987 -447
rect -819 -481 -803 -447
rect -1003 -497 -803 -481
rect -745 -447 -545 -400
rect -745 -481 -729 -447
rect -561 -481 -545 -447
rect -745 -497 -545 -481
rect -487 -447 -287 -400
rect -487 -481 -471 -447
rect -303 -481 -287 -447
rect -487 -497 -287 -481
rect -229 -447 -29 -400
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect -229 -497 -29 -481
rect 29 -447 229 -400
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 29 -497 229 -481
rect 287 -447 487 -400
rect 287 -481 303 -447
rect 471 -481 487 -447
rect 287 -497 487 -481
rect 545 -447 745 -400
rect 545 -481 561 -447
rect 729 -481 745 -447
rect 545 -497 745 -481
rect 803 -447 1003 -400
rect 803 -481 819 -447
rect 987 -481 1003 -447
rect 803 -497 1003 -481
rect 1061 -447 1261 -400
rect 1061 -481 1077 -447
rect 1245 -481 1261 -447
rect 1061 -497 1261 -481
rect 1319 -447 1519 -400
rect 1319 -481 1335 -447
rect 1503 -481 1519 -447
rect 1319 -497 1519 -481
rect 1577 -447 1777 -400
rect 1577 -481 1593 -447
rect 1761 -481 1777 -447
rect 1577 -497 1777 -481
rect 1835 -447 2035 -400
rect 1835 -481 1851 -447
rect 2019 -481 2035 -447
rect 1835 -497 2035 -481
rect 2093 -447 2293 -400
rect 2093 -481 2109 -447
rect 2277 -481 2293 -447
rect 2093 -497 2293 -481
rect 2351 -447 2551 -400
rect 2351 -481 2367 -447
rect 2535 -481 2551 -447
rect 2351 -497 2551 -481
rect 2609 -447 2809 -400
rect 2609 -481 2625 -447
rect 2793 -481 2809 -447
rect 2609 -497 2809 -481
rect 2867 -447 3067 -400
rect 2867 -481 2883 -447
rect 3051 -481 3067 -447
rect 2867 -497 3067 -481
rect 3125 -447 3325 -400
rect 3125 -481 3141 -447
rect 3309 -481 3325 -447
rect 3125 -497 3325 -481
rect 3383 -447 3583 -400
rect 3383 -481 3399 -447
rect 3567 -481 3583 -447
rect 3383 -497 3583 -481
rect 3641 -447 3841 -400
rect 3641 -481 3657 -447
rect 3825 -481 3841 -447
rect 3641 -497 3841 -481
rect 3899 -447 4099 -400
rect 3899 -481 3915 -447
rect 4083 -481 4099 -447
rect 3899 -497 4099 -481
<< polycont >>
rect -4083 447 -3915 481
rect -3825 447 -3657 481
rect -3567 447 -3399 481
rect -3309 447 -3141 481
rect -3051 447 -2883 481
rect -2793 447 -2625 481
rect -2535 447 -2367 481
rect -2277 447 -2109 481
rect -2019 447 -1851 481
rect -1761 447 -1593 481
rect -1503 447 -1335 481
rect -1245 447 -1077 481
rect -987 447 -819 481
rect -729 447 -561 481
rect -471 447 -303 481
rect -213 447 -45 481
rect 45 447 213 481
rect 303 447 471 481
rect 561 447 729 481
rect 819 447 987 481
rect 1077 447 1245 481
rect 1335 447 1503 481
rect 1593 447 1761 481
rect 1851 447 2019 481
rect 2109 447 2277 481
rect 2367 447 2535 481
rect 2625 447 2793 481
rect 2883 447 3051 481
rect 3141 447 3309 481
rect 3399 447 3567 481
rect 3657 447 3825 481
rect 3915 447 4083 481
rect -4083 -481 -3915 -447
rect -3825 -481 -3657 -447
rect -3567 -481 -3399 -447
rect -3309 -481 -3141 -447
rect -3051 -481 -2883 -447
rect -2793 -481 -2625 -447
rect -2535 -481 -2367 -447
rect -2277 -481 -2109 -447
rect -2019 -481 -1851 -447
rect -1761 -481 -1593 -447
rect -1503 -481 -1335 -447
rect -1245 -481 -1077 -447
rect -987 -481 -819 -447
rect -729 -481 -561 -447
rect -471 -481 -303 -447
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect 303 -481 471 -447
rect 561 -481 729 -447
rect 819 -481 987 -447
rect 1077 -481 1245 -447
rect 1335 -481 1503 -447
rect 1593 -481 1761 -447
rect 1851 -481 2019 -447
rect 2109 -481 2277 -447
rect 2367 -481 2535 -447
rect 2625 -481 2793 -447
rect 2883 -481 3051 -447
rect 3141 -481 3309 -447
rect 3399 -481 3567 -447
rect 3657 -481 3825 -447
rect 3915 -481 4083 -447
<< locali >>
rect -4279 585 -4183 619
rect 4183 585 4279 619
rect -4279 523 -4245 585
rect 4245 523 4279 585
rect -4099 447 -4083 481
rect -3915 447 -3899 481
rect -3841 447 -3825 481
rect -3657 447 -3641 481
rect -3583 447 -3567 481
rect -3399 447 -3383 481
rect -3325 447 -3309 481
rect -3141 447 -3125 481
rect -3067 447 -3051 481
rect -2883 447 -2867 481
rect -2809 447 -2793 481
rect -2625 447 -2609 481
rect -2551 447 -2535 481
rect -2367 447 -2351 481
rect -2293 447 -2277 481
rect -2109 447 -2093 481
rect -2035 447 -2019 481
rect -1851 447 -1835 481
rect -1777 447 -1761 481
rect -1593 447 -1577 481
rect -1519 447 -1503 481
rect -1335 447 -1319 481
rect -1261 447 -1245 481
rect -1077 447 -1061 481
rect -1003 447 -987 481
rect -819 447 -803 481
rect -745 447 -729 481
rect -561 447 -545 481
rect -487 447 -471 481
rect -303 447 -287 481
rect -229 447 -213 481
rect -45 447 -29 481
rect 29 447 45 481
rect 213 447 229 481
rect 287 447 303 481
rect 471 447 487 481
rect 545 447 561 481
rect 729 447 745 481
rect 803 447 819 481
rect 987 447 1003 481
rect 1061 447 1077 481
rect 1245 447 1261 481
rect 1319 447 1335 481
rect 1503 447 1519 481
rect 1577 447 1593 481
rect 1761 447 1777 481
rect 1835 447 1851 481
rect 2019 447 2035 481
rect 2093 447 2109 481
rect 2277 447 2293 481
rect 2351 447 2367 481
rect 2535 447 2551 481
rect 2609 447 2625 481
rect 2793 447 2809 481
rect 2867 447 2883 481
rect 3051 447 3067 481
rect 3125 447 3141 481
rect 3309 447 3325 481
rect 3383 447 3399 481
rect 3567 447 3583 481
rect 3641 447 3657 481
rect 3825 447 3841 481
rect 3899 447 3915 481
rect 4083 447 4099 481
rect -4145 388 -4111 404
rect -4145 -404 -4111 -388
rect -3887 388 -3853 404
rect -3887 -404 -3853 -388
rect -3629 388 -3595 404
rect -3629 -404 -3595 -388
rect -3371 388 -3337 404
rect -3371 -404 -3337 -388
rect -3113 388 -3079 404
rect -3113 -404 -3079 -388
rect -2855 388 -2821 404
rect -2855 -404 -2821 -388
rect -2597 388 -2563 404
rect -2597 -404 -2563 -388
rect -2339 388 -2305 404
rect -2339 -404 -2305 -388
rect -2081 388 -2047 404
rect -2081 -404 -2047 -388
rect -1823 388 -1789 404
rect -1823 -404 -1789 -388
rect -1565 388 -1531 404
rect -1565 -404 -1531 -388
rect -1307 388 -1273 404
rect -1307 -404 -1273 -388
rect -1049 388 -1015 404
rect -1049 -404 -1015 -388
rect -791 388 -757 404
rect -791 -404 -757 -388
rect -533 388 -499 404
rect -533 -404 -499 -388
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
rect 499 388 533 404
rect 499 -404 533 -388
rect 757 388 791 404
rect 757 -404 791 -388
rect 1015 388 1049 404
rect 1015 -404 1049 -388
rect 1273 388 1307 404
rect 1273 -404 1307 -388
rect 1531 388 1565 404
rect 1531 -404 1565 -388
rect 1789 388 1823 404
rect 1789 -404 1823 -388
rect 2047 388 2081 404
rect 2047 -404 2081 -388
rect 2305 388 2339 404
rect 2305 -404 2339 -388
rect 2563 388 2597 404
rect 2563 -404 2597 -388
rect 2821 388 2855 404
rect 2821 -404 2855 -388
rect 3079 388 3113 404
rect 3079 -404 3113 -388
rect 3337 388 3371 404
rect 3337 -404 3371 -388
rect 3595 388 3629 404
rect 3595 -404 3629 -388
rect 3853 388 3887 404
rect 3853 -404 3887 -388
rect 4111 388 4145 404
rect 4111 -404 4145 -388
rect -4099 -481 -4083 -447
rect -3915 -481 -3899 -447
rect -3841 -481 -3825 -447
rect -3657 -481 -3641 -447
rect -3583 -481 -3567 -447
rect -3399 -481 -3383 -447
rect -3325 -481 -3309 -447
rect -3141 -481 -3125 -447
rect -3067 -481 -3051 -447
rect -2883 -481 -2867 -447
rect -2809 -481 -2793 -447
rect -2625 -481 -2609 -447
rect -2551 -481 -2535 -447
rect -2367 -481 -2351 -447
rect -2293 -481 -2277 -447
rect -2109 -481 -2093 -447
rect -2035 -481 -2019 -447
rect -1851 -481 -1835 -447
rect -1777 -481 -1761 -447
rect -1593 -481 -1577 -447
rect -1519 -481 -1503 -447
rect -1335 -481 -1319 -447
rect -1261 -481 -1245 -447
rect -1077 -481 -1061 -447
rect -1003 -481 -987 -447
rect -819 -481 -803 -447
rect -745 -481 -729 -447
rect -561 -481 -545 -447
rect -487 -481 -471 -447
rect -303 -481 -287 -447
rect -229 -481 -213 -447
rect -45 -481 -29 -447
rect 29 -481 45 -447
rect 213 -481 229 -447
rect 287 -481 303 -447
rect 471 -481 487 -447
rect 545 -481 561 -447
rect 729 -481 745 -447
rect 803 -481 819 -447
rect 987 -481 1003 -447
rect 1061 -481 1077 -447
rect 1245 -481 1261 -447
rect 1319 -481 1335 -447
rect 1503 -481 1519 -447
rect 1577 -481 1593 -447
rect 1761 -481 1777 -447
rect 1835 -481 1851 -447
rect 2019 -481 2035 -447
rect 2093 -481 2109 -447
rect 2277 -481 2293 -447
rect 2351 -481 2367 -447
rect 2535 -481 2551 -447
rect 2609 -481 2625 -447
rect 2793 -481 2809 -447
rect 2867 -481 2883 -447
rect 3051 -481 3067 -447
rect 3125 -481 3141 -447
rect 3309 -481 3325 -447
rect 3383 -481 3399 -447
rect 3567 -481 3583 -447
rect 3641 -481 3657 -447
rect 3825 -481 3841 -447
rect 3899 -481 3915 -447
rect 4083 -481 4099 -447
rect -4279 -585 -4245 -523
rect 4245 -585 4279 -523
rect -4279 -619 -4183 -585
rect 4183 -619 4279 -585
<< viali >>
rect -4083 447 -3915 481
rect -3825 447 -3657 481
rect -3567 447 -3399 481
rect -3309 447 -3141 481
rect -3051 447 -2883 481
rect -2793 447 -2625 481
rect -2535 447 -2367 481
rect -2277 447 -2109 481
rect -2019 447 -1851 481
rect -1761 447 -1593 481
rect -1503 447 -1335 481
rect -1245 447 -1077 481
rect -987 447 -819 481
rect -729 447 -561 481
rect -471 447 -303 481
rect -213 447 -45 481
rect 45 447 213 481
rect 303 447 471 481
rect 561 447 729 481
rect 819 447 987 481
rect 1077 447 1245 481
rect 1335 447 1503 481
rect 1593 447 1761 481
rect 1851 447 2019 481
rect 2109 447 2277 481
rect 2367 447 2535 481
rect 2625 447 2793 481
rect 2883 447 3051 481
rect 3141 447 3309 481
rect 3399 447 3567 481
rect 3657 447 3825 481
rect 3915 447 4083 481
rect -4145 -388 -4111 388
rect -3887 -388 -3853 388
rect -3629 -388 -3595 388
rect -3371 -388 -3337 388
rect -3113 -388 -3079 388
rect -2855 -388 -2821 388
rect -2597 -388 -2563 388
rect -2339 -388 -2305 388
rect -2081 -388 -2047 388
rect -1823 -388 -1789 388
rect -1565 -388 -1531 388
rect -1307 -388 -1273 388
rect -1049 -388 -1015 388
rect -791 -388 -757 388
rect -533 -388 -499 388
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
rect 499 -388 533 388
rect 757 -388 791 388
rect 1015 -388 1049 388
rect 1273 -388 1307 388
rect 1531 -388 1565 388
rect 1789 -388 1823 388
rect 2047 -388 2081 388
rect 2305 -388 2339 388
rect 2563 -388 2597 388
rect 2821 -388 2855 388
rect 3079 -388 3113 388
rect 3337 -388 3371 388
rect 3595 -388 3629 388
rect 3853 -388 3887 388
rect 4111 -388 4145 388
rect -4083 -481 -3915 -447
rect -3825 -481 -3657 -447
rect -3567 -481 -3399 -447
rect -3309 -481 -3141 -447
rect -3051 -481 -2883 -447
rect -2793 -481 -2625 -447
rect -2535 -481 -2367 -447
rect -2277 -481 -2109 -447
rect -2019 -481 -1851 -447
rect -1761 -481 -1593 -447
rect -1503 -481 -1335 -447
rect -1245 -481 -1077 -447
rect -987 -481 -819 -447
rect -729 -481 -561 -447
rect -471 -481 -303 -447
rect -213 -481 -45 -447
rect 45 -481 213 -447
rect 303 -481 471 -447
rect 561 -481 729 -447
rect 819 -481 987 -447
rect 1077 -481 1245 -447
rect 1335 -481 1503 -447
rect 1593 -481 1761 -447
rect 1851 -481 2019 -447
rect 2109 -481 2277 -447
rect 2367 -481 2535 -447
rect 2625 -481 2793 -447
rect 2883 -481 3051 -447
rect 3141 -481 3309 -447
rect 3399 -481 3567 -447
rect 3657 -481 3825 -447
rect 3915 -481 4083 -447
<< metal1 >>
rect -4095 481 -3903 487
rect -4095 447 -4083 481
rect -3915 447 -3903 481
rect -4095 441 -3903 447
rect -3837 481 -3645 487
rect -3837 447 -3825 481
rect -3657 447 -3645 481
rect -3837 441 -3645 447
rect -3579 481 -3387 487
rect -3579 447 -3567 481
rect -3399 447 -3387 481
rect -3579 441 -3387 447
rect -3321 481 -3129 487
rect -3321 447 -3309 481
rect -3141 447 -3129 481
rect -3321 441 -3129 447
rect -3063 481 -2871 487
rect -3063 447 -3051 481
rect -2883 447 -2871 481
rect -3063 441 -2871 447
rect -2805 481 -2613 487
rect -2805 447 -2793 481
rect -2625 447 -2613 481
rect -2805 441 -2613 447
rect -2547 481 -2355 487
rect -2547 447 -2535 481
rect -2367 447 -2355 481
rect -2547 441 -2355 447
rect -2289 481 -2097 487
rect -2289 447 -2277 481
rect -2109 447 -2097 481
rect -2289 441 -2097 447
rect -2031 481 -1839 487
rect -2031 447 -2019 481
rect -1851 447 -1839 481
rect -2031 441 -1839 447
rect -1773 481 -1581 487
rect -1773 447 -1761 481
rect -1593 447 -1581 481
rect -1773 441 -1581 447
rect -1515 481 -1323 487
rect -1515 447 -1503 481
rect -1335 447 -1323 481
rect -1515 441 -1323 447
rect -1257 481 -1065 487
rect -1257 447 -1245 481
rect -1077 447 -1065 481
rect -1257 441 -1065 447
rect -999 481 -807 487
rect -999 447 -987 481
rect -819 447 -807 481
rect -999 441 -807 447
rect -741 481 -549 487
rect -741 447 -729 481
rect -561 447 -549 481
rect -741 441 -549 447
rect -483 481 -291 487
rect -483 447 -471 481
rect -303 447 -291 481
rect -483 441 -291 447
rect -225 481 -33 487
rect -225 447 -213 481
rect -45 447 -33 481
rect -225 441 -33 447
rect 33 481 225 487
rect 33 447 45 481
rect 213 447 225 481
rect 33 441 225 447
rect 291 481 483 487
rect 291 447 303 481
rect 471 447 483 481
rect 291 441 483 447
rect 549 481 741 487
rect 549 447 561 481
rect 729 447 741 481
rect 549 441 741 447
rect 807 481 999 487
rect 807 447 819 481
rect 987 447 999 481
rect 807 441 999 447
rect 1065 481 1257 487
rect 1065 447 1077 481
rect 1245 447 1257 481
rect 1065 441 1257 447
rect 1323 481 1515 487
rect 1323 447 1335 481
rect 1503 447 1515 481
rect 1323 441 1515 447
rect 1581 481 1773 487
rect 1581 447 1593 481
rect 1761 447 1773 481
rect 1581 441 1773 447
rect 1839 481 2031 487
rect 1839 447 1851 481
rect 2019 447 2031 481
rect 1839 441 2031 447
rect 2097 481 2289 487
rect 2097 447 2109 481
rect 2277 447 2289 481
rect 2097 441 2289 447
rect 2355 481 2547 487
rect 2355 447 2367 481
rect 2535 447 2547 481
rect 2355 441 2547 447
rect 2613 481 2805 487
rect 2613 447 2625 481
rect 2793 447 2805 481
rect 2613 441 2805 447
rect 2871 481 3063 487
rect 2871 447 2883 481
rect 3051 447 3063 481
rect 2871 441 3063 447
rect 3129 481 3321 487
rect 3129 447 3141 481
rect 3309 447 3321 481
rect 3129 441 3321 447
rect 3387 481 3579 487
rect 3387 447 3399 481
rect 3567 447 3579 481
rect 3387 441 3579 447
rect 3645 481 3837 487
rect 3645 447 3657 481
rect 3825 447 3837 481
rect 3645 441 3837 447
rect 3903 481 4095 487
rect 3903 447 3915 481
rect 4083 447 4095 481
rect 3903 441 4095 447
rect -4151 388 -4105 400
rect -4151 -388 -4145 388
rect -4111 -388 -4105 388
rect -4151 -400 -4105 -388
rect -3893 388 -3847 400
rect -3893 -388 -3887 388
rect -3853 -388 -3847 388
rect -3893 -400 -3847 -388
rect -3635 388 -3589 400
rect -3635 -388 -3629 388
rect -3595 -388 -3589 388
rect -3635 -400 -3589 -388
rect -3377 388 -3331 400
rect -3377 -388 -3371 388
rect -3337 -388 -3331 388
rect -3377 -400 -3331 -388
rect -3119 388 -3073 400
rect -3119 -388 -3113 388
rect -3079 -388 -3073 388
rect -3119 -400 -3073 -388
rect -2861 388 -2815 400
rect -2861 -388 -2855 388
rect -2821 -388 -2815 388
rect -2861 -400 -2815 -388
rect -2603 388 -2557 400
rect -2603 -388 -2597 388
rect -2563 -388 -2557 388
rect -2603 -400 -2557 -388
rect -2345 388 -2299 400
rect -2345 -388 -2339 388
rect -2305 -388 -2299 388
rect -2345 -400 -2299 -388
rect -2087 388 -2041 400
rect -2087 -388 -2081 388
rect -2047 -388 -2041 388
rect -2087 -400 -2041 -388
rect -1829 388 -1783 400
rect -1829 -388 -1823 388
rect -1789 -388 -1783 388
rect -1829 -400 -1783 -388
rect -1571 388 -1525 400
rect -1571 -388 -1565 388
rect -1531 -388 -1525 388
rect -1571 -400 -1525 -388
rect -1313 388 -1267 400
rect -1313 -388 -1307 388
rect -1273 -388 -1267 388
rect -1313 -400 -1267 -388
rect -1055 388 -1009 400
rect -1055 -388 -1049 388
rect -1015 -388 -1009 388
rect -1055 -400 -1009 -388
rect -797 388 -751 400
rect -797 -388 -791 388
rect -757 -388 -751 388
rect -797 -400 -751 -388
rect -539 388 -493 400
rect -539 -388 -533 388
rect -499 -388 -493 388
rect -539 -400 -493 -388
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
rect 493 388 539 400
rect 493 -388 499 388
rect 533 -388 539 388
rect 493 -400 539 -388
rect 751 388 797 400
rect 751 -388 757 388
rect 791 -388 797 388
rect 751 -400 797 -388
rect 1009 388 1055 400
rect 1009 -388 1015 388
rect 1049 -388 1055 388
rect 1009 -400 1055 -388
rect 1267 388 1313 400
rect 1267 -388 1273 388
rect 1307 -388 1313 388
rect 1267 -400 1313 -388
rect 1525 388 1571 400
rect 1525 -388 1531 388
rect 1565 -388 1571 388
rect 1525 -400 1571 -388
rect 1783 388 1829 400
rect 1783 -388 1789 388
rect 1823 -388 1829 388
rect 1783 -400 1829 -388
rect 2041 388 2087 400
rect 2041 -388 2047 388
rect 2081 -388 2087 388
rect 2041 -400 2087 -388
rect 2299 388 2345 400
rect 2299 -388 2305 388
rect 2339 -388 2345 388
rect 2299 -400 2345 -388
rect 2557 388 2603 400
rect 2557 -388 2563 388
rect 2597 -388 2603 388
rect 2557 -400 2603 -388
rect 2815 388 2861 400
rect 2815 -388 2821 388
rect 2855 -388 2861 388
rect 2815 -400 2861 -388
rect 3073 388 3119 400
rect 3073 -388 3079 388
rect 3113 -388 3119 388
rect 3073 -400 3119 -388
rect 3331 388 3377 400
rect 3331 -388 3337 388
rect 3371 -388 3377 388
rect 3331 -400 3377 -388
rect 3589 388 3635 400
rect 3589 -388 3595 388
rect 3629 -388 3635 388
rect 3589 -400 3635 -388
rect 3847 388 3893 400
rect 3847 -388 3853 388
rect 3887 -388 3893 388
rect 3847 -400 3893 -388
rect 4105 388 4151 400
rect 4105 -388 4111 388
rect 4145 -388 4151 388
rect 4105 -400 4151 -388
rect -4095 -447 -3903 -441
rect -4095 -481 -4083 -447
rect -3915 -481 -3903 -447
rect -4095 -487 -3903 -481
rect -3837 -447 -3645 -441
rect -3837 -481 -3825 -447
rect -3657 -481 -3645 -447
rect -3837 -487 -3645 -481
rect -3579 -447 -3387 -441
rect -3579 -481 -3567 -447
rect -3399 -481 -3387 -447
rect -3579 -487 -3387 -481
rect -3321 -447 -3129 -441
rect -3321 -481 -3309 -447
rect -3141 -481 -3129 -447
rect -3321 -487 -3129 -481
rect -3063 -447 -2871 -441
rect -3063 -481 -3051 -447
rect -2883 -481 -2871 -447
rect -3063 -487 -2871 -481
rect -2805 -447 -2613 -441
rect -2805 -481 -2793 -447
rect -2625 -481 -2613 -447
rect -2805 -487 -2613 -481
rect -2547 -447 -2355 -441
rect -2547 -481 -2535 -447
rect -2367 -481 -2355 -447
rect -2547 -487 -2355 -481
rect -2289 -447 -2097 -441
rect -2289 -481 -2277 -447
rect -2109 -481 -2097 -447
rect -2289 -487 -2097 -481
rect -2031 -447 -1839 -441
rect -2031 -481 -2019 -447
rect -1851 -481 -1839 -447
rect -2031 -487 -1839 -481
rect -1773 -447 -1581 -441
rect -1773 -481 -1761 -447
rect -1593 -481 -1581 -447
rect -1773 -487 -1581 -481
rect -1515 -447 -1323 -441
rect -1515 -481 -1503 -447
rect -1335 -481 -1323 -447
rect -1515 -487 -1323 -481
rect -1257 -447 -1065 -441
rect -1257 -481 -1245 -447
rect -1077 -481 -1065 -447
rect -1257 -487 -1065 -481
rect -999 -447 -807 -441
rect -999 -481 -987 -447
rect -819 -481 -807 -447
rect -999 -487 -807 -481
rect -741 -447 -549 -441
rect -741 -481 -729 -447
rect -561 -481 -549 -447
rect -741 -487 -549 -481
rect -483 -447 -291 -441
rect -483 -481 -471 -447
rect -303 -481 -291 -447
rect -483 -487 -291 -481
rect -225 -447 -33 -441
rect -225 -481 -213 -447
rect -45 -481 -33 -447
rect -225 -487 -33 -481
rect 33 -447 225 -441
rect 33 -481 45 -447
rect 213 -481 225 -447
rect 33 -487 225 -481
rect 291 -447 483 -441
rect 291 -481 303 -447
rect 471 -481 483 -447
rect 291 -487 483 -481
rect 549 -447 741 -441
rect 549 -481 561 -447
rect 729 -481 741 -447
rect 549 -487 741 -481
rect 807 -447 999 -441
rect 807 -481 819 -447
rect 987 -481 999 -447
rect 807 -487 999 -481
rect 1065 -447 1257 -441
rect 1065 -481 1077 -447
rect 1245 -481 1257 -447
rect 1065 -487 1257 -481
rect 1323 -447 1515 -441
rect 1323 -481 1335 -447
rect 1503 -481 1515 -447
rect 1323 -487 1515 -481
rect 1581 -447 1773 -441
rect 1581 -481 1593 -447
rect 1761 -481 1773 -447
rect 1581 -487 1773 -481
rect 1839 -447 2031 -441
rect 1839 -481 1851 -447
rect 2019 -481 2031 -447
rect 1839 -487 2031 -481
rect 2097 -447 2289 -441
rect 2097 -481 2109 -447
rect 2277 -481 2289 -447
rect 2097 -487 2289 -481
rect 2355 -447 2547 -441
rect 2355 -481 2367 -447
rect 2535 -481 2547 -447
rect 2355 -487 2547 -481
rect 2613 -447 2805 -441
rect 2613 -481 2625 -447
rect 2793 -481 2805 -447
rect 2613 -487 2805 -481
rect 2871 -447 3063 -441
rect 2871 -481 2883 -447
rect 3051 -481 3063 -447
rect 2871 -487 3063 -481
rect 3129 -447 3321 -441
rect 3129 -481 3141 -447
rect 3309 -481 3321 -447
rect 3129 -487 3321 -481
rect 3387 -447 3579 -441
rect 3387 -481 3399 -447
rect 3567 -481 3579 -447
rect 3387 -487 3579 -481
rect 3645 -447 3837 -441
rect 3645 -481 3657 -447
rect 3825 -481 3837 -447
rect 3645 -487 3837 -481
rect 3903 -447 4095 -441
rect 3903 -481 3915 -447
rect 4083 -481 4095 -447
rect 3903 -487 4095 -481
<< properties >>
string FIXED_BBOX -4262 -602 4262 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 32 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
timestamp 1713232886
<< pwell >>
rect -938 -229 938 229
<< mvnmos >>
rect -824 -100 -724 100
rect -695 -100 -595 100
rect -566 -100 -466 100
rect -437 -100 -337 100
rect -308 -100 -208 100
rect -179 -100 -79 100
rect -50 -100 50 100
rect 79 -100 179 100
rect 208 -100 308 100
rect 337 -100 437 100
rect 466 -100 566 100
rect 595 -100 695 100
rect 724 -100 824 100
<< mvndiff >>
rect -853 94 -824 100
rect -853 -94 -847 94
rect -830 -94 -824 94
rect -853 -100 -824 -94
rect -724 94 -695 100
rect -724 -94 -718 94
rect -701 -94 -695 94
rect -724 -100 -695 -94
rect -595 94 -566 100
rect -595 -94 -589 94
rect -572 -94 -566 94
rect -595 -100 -566 -94
rect -466 94 -437 100
rect -466 -94 -460 94
rect -443 -94 -437 94
rect -466 -100 -437 -94
rect -337 94 -308 100
rect -337 -94 -331 94
rect -314 -94 -308 94
rect -337 -100 -308 -94
rect -208 94 -179 100
rect -208 -94 -202 94
rect -185 -94 -179 94
rect -208 -100 -179 -94
rect -79 94 -50 100
rect -79 -94 -73 94
rect -56 -94 -50 94
rect -79 -100 -50 -94
rect 50 94 79 100
rect 50 -94 56 94
rect 73 -94 79 94
rect 50 -100 79 -94
rect 179 94 208 100
rect 179 -94 185 94
rect 202 -94 208 94
rect 179 -100 208 -94
rect 308 94 337 100
rect 308 -94 314 94
rect 331 -94 337 94
rect 308 -100 337 -94
rect 437 94 466 100
rect 437 -94 443 94
rect 460 -94 466 94
rect 437 -100 466 -94
rect 566 94 595 100
rect 566 -94 572 94
rect 589 -94 595 94
rect 566 -100 595 -94
rect 695 94 724 100
rect 695 -94 701 94
rect 718 -94 724 94
rect 695 -100 724 -94
rect 824 94 853 100
rect 824 -94 830 94
rect 847 -94 853 94
rect 824 -100 853 -94
<< mvndiffc >>
rect -847 -94 -830 94
rect -718 -94 -701 94
rect -589 -94 -572 94
rect -460 -94 -443 94
rect -331 -94 -314 94
rect -202 -94 -185 94
rect -73 -94 -56 94
rect 56 -94 73 94
rect 185 -94 202 94
rect 314 -94 331 94
rect 443 -94 460 94
rect 572 -94 589 94
rect 701 -94 718 94
rect 830 -94 847 94
<< mvpsubdiff >>
rect -920 205 920 211
rect -920 188 -866 205
rect 866 188 920 205
rect -920 182 920 188
rect -920 157 -891 182
rect -920 -157 -914 157
rect -897 -157 -891 157
rect 891 157 920 182
rect -920 -182 -891 -157
rect 891 -157 897 157
rect 914 -157 920 157
rect 891 -182 920 -157
rect -920 -188 920 -182
rect -920 -205 -866 -188
rect 866 -205 920 -188
rect -920 -211 920 -205
<< mvpsubdiffcont >>
rect -866 188 866 205
rect -914 -157 -897 157
rect 897 -157 914 157
rect -866 -205 866 -188
<< poly >>
rect -824 136 -724 144
rect -824 119 -816 136
rect -732 119 -724 136
rect -824 100 -724 119
rect -695 136 -595 144
rect -695 119 -687 136
rect -603 119 -595 136
rect -695 100 -595 119
rect -566 136 -466 144
rect -566 119 -558 136
rect -474 119 -466 136
rect -566 100 -466 119
rect -437 136 -337 144
rect -437 119 -429 136
rect -345 119 -337 136
rect -437 100 -337 119
rect -308 136 -208 144
rect -308 119 -300 136
rect -216 119 -208 136
rect -308 100 -208 119
rect -179 136 -79 144
rect -179 119 -171 136
rect -87 119 -79 136
rect -179 100 -79 119
rect -50 136 50 144
rect -50 119 -42 136
rect 42 119 50 136
rect -50 100 50 119
rect 79 136 179 144
rect 79 119 87 136
rect 171 119 179 136
rect 79 100 179 119
rect 208 136 308 144
rect 208 119 216 136
rect 300 119 308 136
rect 208 100 308 119
rect 337 136 437 144
rect 337 119 345 136
rect 429 119 437 136
rect 337 100 437 119
rect 466 136 566 144
rect 466 119 474 136
rect 558 119 566 136
rect 466 100 566 119
rect 595 136 695 144
rect 595 119 603 136
rect 687 119 695 136
rect 595 100 695 119
rect 724 136 824 144
rect 724 119 732 136
rect 816 119 824 136
rect 724 100 824 119
rect -824 -119 -724 -100
rect -824 -136 -816 -119
rect -732 -136 -724 -119
rect -824 -144 -724 -136
rect -695 -119 -595 -100
rect -695 -136 -687 -119
rect -603 -136 -595 -119
rect -695 -144 -595 -136
rect -566 -119 -466 -100
rect -566 -136 -558 -119
rect -474 -136 -466 -119
rect -566 -144 -466 -136
rect -437 -119 -337 -100
rect -437 -136 -429 -119
rect -345 -136 -337 -119
rect -437 -144 -337 -136
rect -308 -119 -208 -100
rect -308 -136 -300 -119
rect -216 -136 -208 -119
rect -308 -144 -208 -136
rect -179 -119 -79 -100
rect -179 -136 -171 -119
rect -87 -136 -79 -119
rect -179 -144 -79 -136
rect -50 -119 50 -100
rect -50 -136 -42 -119
rect 42 -136 50 -119
rect -50 -144 50 -136
rect 79 -119 179 -100
rect 79 -136 87 -119
rect 171 -136 179 -119
rect 79 -144 179 -136
rect 208 -119 308 -100
rect 208 -136 216 -119
rect 300 -136 308 -119
rect 208 -144 308 -136
rect 337 -119 437 -100
rect 337 -136 345 -119
rect 429 -136 437 -119
rect 337 -144 437 -136
rect 466 -119 566 -100
rect 466 -136 474 -119
rect 558 -136 566 -119
rect 466 -144 566 -136
rect 595 -119 695 -100
rect 595 -136 603 -119
rect 687 -136 695 -119
rect 595 -144 695 -136
rect 724 -119 824 -100
rect 724 -136 732 -119
rect 816 -136 824 -119
rect 724 -144 824 -136
<< polycont >>
rect -816 119 -732 136
rect -687 119 -603 136
rect -558 119 -474 136
rect -429 119 -345 136
rect -300 119 -216 136
rect -171 119 -87 136
rect -42 119 42 136
rect 87 119 171 136
rect 216 119 300 136
rect 345 119 429 136
rect 474 119 558 136
rect 603 119 687 136
rect 732 119 816 136
rect -816 -136 -732 -119
rect -687 -136 -603 -119
rect -558 -136 -474 -119
rect -429 -136 -345 -119
rect -300 -136 -216 -119
rect -171 -136 -87 -119
rect -42 -136 42 -119
rect 87 -136 171 -119
rect 216 -136 300 -119
rect 345 -136 429 -119
rect 474 -136 558 -119
rect 603 -136 687 -119
rect 732 -136 816 -119
<< locali >>
rect -914 188 -866 205
rect 866 188 914 205
rect -914 157 -897 188
rect 897 157 914 188
rect -824 119 -816 136
rect -732 119 -724 136
rect -695 119 -687 136
rect -603 119 -595 136
rect -566 119 -558 136
rect -474 119 -466 136
rect -437 119 -429 136
rect -345 119 -337 136
rect -308 119 -300 136
rect -216 119 -208 136
rect -179 119 -171 136
rect -87 119 -79 136
rect -50 119 -42 136
rect 42 119 50 136
rect 79 119 87 136
rect 171 119 179 136
rect 208 119 216 136
rect 300 119 308 136
rect 337 119 345 136
rect 429 119 437 136
rect 466 119 474 136
rect 558 119 566 136
rect 595 119 603 136
rect 687 119 695 136
rect 724 119 732 136
rect 816 119 824 136
rect -847 94 -830 102
rect -847 -102 -830 -94
rect -718 94 -701 102
rect -718 -102 -701 -94
rect -589 94 -572 102
rect -589 -102 -572 -94
rect -460 94 -443 102
rect -460 -102 -443 -94
rect -331 94 -314 102
rect -331 -102 -314 -94
rect -202 94 -185 102
rect -202 -102 -185 -94
rect -73 94 -56 102
rect -73 -102 -56 -94
rect 56 94 73 102
rect 56 -102 73 -94
rect 185 94 202 102
rect 185 -102 202 -94
rect 314 94 331 102
rect 314 -102 331 -94
rect 443 94 460 102
rect 443 -102 460 -94
rect 572 94 589 102
rect 572 -102 589 -94
rect 701 94 718 102
rect 701 -102 718 -94
rect 830 94 847 102
rect 830 -102 847 -94
rect -824 -136 -816 -119
rect -732 -136 -724 -119
rect -695 -136 -687 -119
rect -603 -136 -595 -119
rect -566 -136 -558 -119
rect -474 -136 -466 -119
rect -437 -136 -429 -119
rect -345 -136 -337 -119
rect -308 -136 -300 -119
rect -216 -136 -208 -119
rect -179 -136 -171 -119
rect -87 -136 -79 -119
rect -50 -136 -42 -119
rect 42 -136 50 -119
rect 79 -136 87 -119
rect 171 -136 179 -119
rect 208 -136 216 -119
rect 300 -136 308 -119
rect 337 -136 345 -119
rect 429 -136 437 -119
rect 466 -136 474 -119
rect 558 -136 566 -119
rect 595 -136 603 -119
rect 687 -136 695 -119
rect 724 -136 732 -119
rect 816 -136 824 -119
rect -914 -188 -897 -157
rect 897 -188 914 -157
rect -914 -205 -866 -188
rect 866 -205 914 -188
<< viali >>
rect -816 119 -732 136
rect -687 119 -603 136
rect -558 119 -474 136
rect -429 119 -345 136
rect -300 119 -216 136
rect -171 119 -87 136
rect -42 119 42 136
rect 87 119 171 136
rect 216 119 300 136
rect 345 119 429 136
rect 474 119 558 136
rect 603 119 687 136
rect 732 119 816 136
rect -847 -94 -830 94
rect -718 -94 -701 94
rect -589 -94 -572 94
rect -460 -94 -443 94
rect -331 -94 -314 94
rect -202 -94 -185 94
rect -73 -94 -56 94
rect 56 -94 73 94
rect 185 -94 202 94
rect 314 -94 331 94
rect 443 -94 460 94
rect 572 -94 589 94
rect 701 -94 718 94
rect 830 -94 847 94
rect -816 -136 -732 -119
rect -687 -136 -603 -119
rect -558 -136 -474 -119
rect -429 -136 -345 -119
rect -300 -136 -216 -119
rect -171 -136 -87 -119
rect -42 -136 42 -119
rect 87 -136 171 -119
rect 216 -136 300 -119
rect 345 -136 429 -119
rect 474 -136 558 -119
rect 603 -136 687 -119
rect 732 -136 816 -119
<< metal1 >>
rect -822 136 -726 139
rect -822 119 -816 136
rect -732 119 -726 136
rect -822 116 -726 119
rect -693 136 -597 139
rect -693 119 -687 136
rect -603 119 -597 136
rect -693 116 -597 119
rect -564 136 -468 139
rect -564 119 -558 136
rect -474 119 -468 136
rect -564 116 -468 119
rect -435 136 -339 139
rect -435 119 -429 136
rect -345 119 -339 136
rect -435 116 -339 119
rect -306 136 -210 139
rect -306 119 -300 136
rect -216 119 -210 136
rect -306 116 -210 119
rect -177 136 -81 139
rect -177 119 -171 136
rect -87 119 -81 136
rect -177 116 -81 119
rect -48 136 48 139
rect -48 119 -42 136
rect 42 119 48 136
rect -48 116 48 119
rect 81 136 177 139
rect 81 119 87 136
rect 171 119 177 136
rect 81 116 177 119
rect 210 136 306 139
rect 210 119 216 136
rect 300 119 306 136
rect 210 116 306 119
rect 339 136 435 139
rect 339 119 345 136
rect 429 119 435 136
rect 339 116 435 119
rect 468 136 564 139
rect 468 119 474 136
rect 558 119 564 136
rect 468 116 564 119
rect 597 136 693 139
rect 597 119 603 136
rect 687 119 693 136
rect 597 116 693 119
rect 726 136 822 139
rect 726 119 732 136
rect 816 119 822 136
rect 726 116 822 119
rect -850 94 -827 100
rect -850 -94 -847 94
rect -830 -94 -827 94
rect -850 -100 -827 -94
rect -721 94 -698 100
rect -721 -94 -718 94
rect -701 -94 -698 94
rect -721 -100 -698 -94
rect -592 94 -569 100
rect -592 -94 -589 94
rect -572 -94 -569 94
rect -592 -100 -569 -94
rect -463 94 -440 100
rect -463 -94 -460 94
rect -443 -94 -440 94
rect -463 -100 -440 -94
rect -334 94 -311 100
rect -334 -94 -331 94
rect -314 -94 -311 94
rect -334 -100 -311 -94
rect -205 94 -182 100
rect -205 -94 -202 94
rect -185 -94 -182 94
rect -205 -100 -182 -94
rect -76 94 -53 100
rect -76 -94 -73 94
rect -56 -94 -53 94
rect -76 -100 -53 -94
rect 53 94 76 100
rect 53 -94 56 94
rect 73 -94 76 94
rect 53 -100 76 -94
rect 182 94 205 100
rect 182 -94 185 94
rect 202 -94 205 94
rect 182 -100 205 -94
rect 311 94 334 100
rect 311 -94 314 94
rect 331 -94 334 94
rect 311 -100 334 -94
rect 440 94 463 100
rect 440 -94 443 94
rect 460 -94 463 94
rect 440 -100 463 -94
rect 569 94 592 100
rect 569 -94 572 94
rect 589 -94 592 94
rect 569 -100 592 -94
rect 698 94 721 100
rect 698 -94 701 94
rect 718 -94 721 94
rect 698 -100 721 -94
rect 827 94 850 100
rect 827 -94 830 94
rect 847 -94 850 94
rect 827 -100 850 -94
rect -822 -119 -726 -116
rect -822 -136 -816 -119
rect -732 -136 -726 -119
rect -822 -139 -726 -136
rect -693 -119 -597 -116
rect -693 -136 -687 -119
rect -603 -136 -597 -119
rect -693 -139 -597 -136
rect -564 -119 -468 -116
rect -564 -136 -558 -119
rect -474 -136 -468 -119
rect -564 -139 -468 -136
rect -435 -119 -339 -116
rect -435 -136 -429 -119
rect -345 -136 -339 -119
rect -435 -139 -339 -136
rect -306 -119 -210 -116
rect -306 -136 -300 -119
rect -216 -136 -210 -119
rect -306 -139 -210 -136
rect -177 -119 -81 -116
rect -177 -136 -171 -119
rect -87 -136 -81 -119
rect -177 -139 -81 -136
rect -48 -119 48 -116
rect -48 -136 -42 -119
rect 42 -136 48 -119
rect -48 -139 48 -136
rect 81 -119 177 -116
rect 81 -136 87 -119
rect 171 -136 177 -119
rect 81 -139 177 -136
rect 210 -119 306 -116
rect 210 -136 216 -119
rect 300 -136 306 -119
rect 210 -139 306 -136
rect 339 -119 435 -116
rect 339 -136 345 -119
rect 429 -136 435 -119
rect 339 -139 435 -136
rect 468 -119 564 -116
rect 468 -136 474 -119
rect 558 -136 564 -119
rect 468 -139 564 -136
rect 597 -119 693 -116
rect 597 -136 603 -119
rect 687 -136 693 -119
rect 597 -139 693 -136
rect 726 -119 822 -116
rect 726 -136 732 -119
rect 816 -136 822 -119
rect 726 -139 822 -136
<< properties >>
string FIXED_BBOX -905 -196 905 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713400206
<< nwell >>
rect -2551 -1897 2551 1897
<< mvpmos >>
rect -2293 -1600 -2093 1600
rect -2035 -1600 -1835 1600
rect -1777 -1600 -1577 1600
rect -1519 -1600 -1319 1600
rect -1261 -1600 -1061 1600
rect -1003 -1600 -803 1600
rect -745 -1600 -545 1600
rect -487 -1600 -287 1600
rect -229 -1600 -29 1600
rect 29 -1600 229 1600
rect 287 -1600 487 1600
rect 545 -1600 745 1600
rect 803 -1600 1003 1600
rect 1061 -1600 1261 1600
rect 1319 -1600 1519 1600
rect 1577 -1600 1777 1600
rect 1835 -1600 2035 1600
rect 2093 -1600 2293 1600
<< mvpdiff >>
rect -2351 1588 -2293 1600
rect -2351 -1588 -2339 1588
rect -2305 -1588 -2293 1588
rect -2351 -1600 -2293 -1588
rect -2093 1588 -2035 1600
rect -2093 -1588 -2081 1588
rect -2047 -1588 -2035 1588
rect -2093 -1600 -2035 -1588
rect -1835 1588 -1777 1600
rect -1835 -1588 -1823 1588
rect -1789 -1588 -1777 1588
rect -1835 -1600 -1777 -1588
rect -1577 1588 -1519 1600
rect -1577 -1588 -1565 1588
rect -1531 -1588 -1519 1588
rect -1577 -1600 -1519 -1588
rect -1319 1588 -1261 1600
rect -1319 -1588 -1307 1588
rect -1273 -1588 -1261 1588
rect -1319 -1600 -1261 -1588
rect -1061 1588 -1003 1600
rect -1061 -1588 -1049 1588
rect -1015 -1588 -1003 1588
rect -1061 -1600 -1003 -1588
rect -803 1588 -745 1600
rect -803 -1588 -791 1588
rect -757 -1588 -745 1588
rect -803 -1600 -745 -1588
rect -545 1588 -487 1600
rect -545 -1588 -533 1588
rect -499 -1588 -487 1588
rect -545 -1600 -487 -1588
rect -287 1588 -229 1600
rect -287 -1588 -275 1588
rect -241 -1588 -229 1588
rect -287 -1600 -229 -1588
rect -29 1588 29 1600
rect -29 -1588 -17 1588
rect 17 -1588 29 1588
rect -29 -1600 29 -1588
rect 229 1588 287 1600
rect 229 -1588 241 1588
rect 275 -1588 287 1588
rect 229 -1600 287 -1588
rect 487 1588 545 1600
rect 487 -1588 499 1588
rect 533 -1588 545 1588
rect 487 -1600 545 -1588
rect 745 1588 803 1600
rect 745 -1588 757 1588
rect 791 -1588 803 1588
rect 745 -1600 803 -1588
rect 1003 1588 1061 1600
rect 1003 -1588 1015 1588
rect 1049 -1588 1061 1588
rect 1003 -1600 1061 -1588
rect 1261 1588 1319 1600
rect 1261 -1588 1273 1588
rect 1307 -1588 1319 1588
rect 1261 -1600 1319 -1588
rect 1519 1588 1577 1600
rect 1519 -1588 1531 1588
rect 1565 -1588 1577 1588
rect 1519 -1600 1577 -1588
rect 1777 1588 1835 1600
rect 1777 -1588 1789 1588
rect 1823 -1588 1835 1588
rect 1777 -1600 1835 -1588
rect 2035 1588 2093 1600
rect 2035 -1588 2047 1588
rect 2081 -1588 2093 1588
rect 2035 -1600 2093 -1588
rect 2293 1588 2351 1600
rect 2293 -1588 2305 1588
rect 2339 -1588 2351 1588
rect 2293 -1600 2351 -1588
<< mvpdiffc >>
rect -2339 -1588 -2305 1588
rect -2081 -1588 -2047 1588
rect -1823 -1588 -1789 1588
rect -1565 -1588 -1531 1588
rect -1307 -1588 -1273 1588
rect -1049 -1588 -1015 1588
rect -791 -1588 -757 1588
rect -533 -1588 -499 1588
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
rect 499 -1588 533 1588
rect 757 -1588 791 1588
rect 1015 -1588 1049 1588
rect 1273 -1588 1307 1588
rect 1531 -1588 1565 1588
rect 1789 -1588 1823 1588
rect 2047 -1588 2081 1588
rect 2305 -1588 2339 1588
<< mvnsubdiff >>
rect -2485 1819 2485 1831
rect -2485 1785 -2377 1819
rect 2377 1785 2485 1819
rect -2485 1773 2485 1785
rect -2485 1723 -2427 1773
rect -2485 -1723 -2473 1723
rect -2439 -1723 -2427 1723
rect 2427 1723 2485 1773
rect -2485 -1773 -2427 -1723
rect 2427 -1723 2439 1723
rect 2473 -1723 2485 1723
rect 2427 -1773 2485 -1723
rect -2485 -1785 2485 -1773
rect -2485 -1819 -2377 -1785
rect 2377 -1819 2485 -1785
rect -2485 -1831 2485 -1819
<< mvnsubdiffcont >>
rect -2377 1785 2377 1819
rect -2473 -1723 -2439 1723
rect 2439 -1723 2473 1723
rect -2377 -1819 2377 -1785
<< poly >>
rect -2259 1681 -2127 1697
rect -2259 1664 -2243 1681
rect -2293 1647 -2243 1664
rect -2143 1664 -2127 1681
rect -2001 1681 -1869 1697
rect -2001 1664 -1985 1681
rect -2143 1647 -2093 1664
rect -2293 1600 -2093 1647
rect -2035 1647 -1985 1664
rect -1885 1664 -1869 1681
rect -1743 1681 -1611 1697
rect -1743 1664 -1727 1681
rect -1885 1647 -1835 1664
rect -2035 1600 -1835 1647
rect -1777 1647 -1727 1664
rect -1627 1664 -1611 1681
rect -1485 1681 -1353 1697
rect -1485 1664 -1469 1681
rect -1627 1647 -1577 1664
rect -1777 1600 -1577 1647
rect -1519 1647 -1469 1664
rect -1369 1664 -1353 1681
rect -1227 1681 -1095 1697
rect -1227 1664 -1211 1681
rect -1369 1647 -1319 1664
rect -1519 1600 -1319 1647
rect -1261 1647 -1211 1664
rect -1111 1664 -1095 1681
rect -969 1681 -837 1697
rect -969 1664 -953 1681
rect -1111 1647 -1061 1664
rect -1261 1600 -1061 1647
rect -1003 1647 -953 1664
rect -853 1664 -837 1681
rect -711 1681 -579 1697
rect -711 1664 -695 1681
rect -853 1647 -803 1664
rect -1003 1600 -803 1647
rect -745 1647 -695 1664
rect -595 1664 -579 1681
rect -453 1681 -321 1697
rect -453 1664 -437 1681
rect -595 1647 -545 1664
rect -745 1600 -545 1647
rect -487 1647 -437 1664
rect -337 1664 -321 1681
rect -195 1681 -63 1697
rect -195 1664 -179 1681
rect -337 1647 -287 1664
rect -487 1600 -287 1647
rect -229 1647 -179 1664
rect -79 1664 -63 1681
rect 63 1681 195 1697
rect 63 1664 79 1681
rect -79 1647 -29 1664
rect -229 1600 -29 1647
rect 29 1647 79 1664
rect 179 1664 195 1681
rect 321 1681 453 1697
rect 321 1664 337 1681
rect 179 1647 229 1664
rect 29 1600 229 1647
rect 287 1647 337 1664
rect 437 1664 453 1681
rect 579 1681 711 1697
rect 579 1664 595 1681
rect 437 1647 487 1664
rect 287 1600 487 1647
rect 545 1647 595 1664
rect 695 1664 711 1681
rect 837 1681 969 1697
rect 837 1664 853 1681
rect 695 1647 745 1664
rect 545 1600 745 1647
rect 803 1647 853 1664
rect 953 1664 969 1681
rect 1095 1681 1227 1697
rect 1095 1664 1111 1681
rect 953 1647 1003 1664
rect 803 1600 1003 1647
rect 1061 1647 1111 1664
rect 1211 1664 1227 1681
rect 1353 1681 1485 1697
rect 1353 1664 1369 1681
rect 1211 1647 1261 1664
rect 1061 1600 1261 1647
rect 1319 1647 1369 1664
rect 1469 1664 1485 1681
rect 1611 1681 1743 1697
rect 1611 1664 1627 1681
rect 1469 1647 1519 1664
rect 1319 1600 1519 1647
rect 1577 1647 1627 1664
rect 1727 1664 1743 1681
rect 1869 1681 2001 1697
rect 1869 1664 1885 1681
rect 1727 1647 1777 1664
rect 1577 1600 1777 1647
rect 1835 1647 1885 1664
rect 1985 1664 2001 1681
rect 2127 1681 2259 1697
rect 2127 1664 2143 1681
rect 1985 1647 2035 1664
rect 1835 1600 2035 1647
rect 2093 1647 2143 1664
rect 2243 1664 2259 1681
rect 2243 1647 2293 1664
rect 2093 1600 2293 1647
rect -2293 -1647 -2093 -1600
rect -2293 -1664 -2243 -1647
rect -2259 -1681 -2243 -1664
rect -2143 -1664 -2093 -1647
rect -2035 -1647 -1835 -1600
rect -2035 -1664 -1985 -1647
rect -2143 -1681 -2127 -1664
rect -2259 -1697 -2127 -1681
rect -2001 -1681 -1985 -1664
rect -1885 -1664 -1835 -1647
rect -1777 -1647 -1577 -1600
rect -1777 -1664 -1727 -1647
rect -1885 -1681 -1869 -1664
rect -2001 -1697 -1869 -1681
rect -1743 -1681 -1727 -1664
rect -1627 -1664 -1577 -1647
rect -1519 -1647 -1319 -1600
rect -1519 -1664 -1469 -1647
rect -1627 -1681 -1611 -1664
rect -1743 -1697 -1611 -1681
rect -1485 -1681 -1469 -1664
rect -1369 -1664 -1319 -1647
rect -1261 -1647 -1061 -1600
rect -1261 -1664 -1211 -1647
rect -1369 -1681 -1353 -1664
rect -1485 -1697 -1353 -1681
rect -1227 -1681 -1211 -1664
rect -1111 -1664 -1061 -1647
rect -1003 -1647 -803 -1600
rect -1003 -1664 -953 -1647
rect -1111 -1681 -1095 -1664
rect -1227 -1697 -1095 -1681
rect -969 -1681 -953 -1664
rect -853 -1664 -803 -1647
rect -745 -1647 -545 -1600
rect -745 -1664 -695 -1647
rect -853 -1681 -837 -1664
rect -969 -1697 -837 -1681
rect -711 -1681 -695 -1664
rect -595 -1664 -545 -1647
rect -487 -1647 -287 -1600
rect -487 -1664 -437 -1647
rect -595 -1681 -579 -1664
rect -711 -1697 -579 -1681
rect -453 -1681 -437 -1664
rect -337 -1664 -287 -1647
rect -229 -1647 -29 -1600
rect -229 -1664 -179 -1647
rect -337 -1681 -321 -1664
rect -453 -1697 -321 -1681
rect -195 -1681 -179 -1664
rect -79 -1664 -29 -1647
rect 29 -1647 229 -1600
rect 29 -1664 79 -1647
rect -79 -1681 -63 -1664
rect -195 -1697 -63 -1681
rect 63 -1681 79 -1664
rect 179 -1664 229 -1647
rect 287 -1647 487 -1600
rect 287 -1664 337 -1647
rect 179 -1681 195 -1664
rect 63 -1697 195 -1681
rect 321 -1681 337 -1664
rect 437 -1664 487 -1647
rect 545 -1647 745 -1600
rect 545 -1664 595 -1647
rect 437 -1681 453 -1664
rect 321 -1697 453 -1681
rect 579 -1681 595 -1664
rect 695 -1664 745 -1647
rect 803 -1647 1003 -1600
rect 803 -1664 853 -1647
rect 695 -1681 711 -1664
rect 579 -1697 711 -1681
rect 837 -1681 853 -1664
rect 953 -1664 1003 -1647
rect 1061 -1647 1261 -1600
rect 1061 -1664 1111 -1647
rect 953 -1681 969 -1664
rect 837 -1697 969 -1681
rect 1095 -1681 1111 -1664
rect 1211 -1664 1261 -1647
rect 1319 -1647 1519 -1600
rect 1319 -1664 1369 -1647
rect 1211 -1681 1227 -1664
rect 1095 -1697 1227 -1681
rect 1353 -1681 1369 -1664
rect 1469 -1664 1519 -1647
rect 1577 -1647 1777 -1600
rect 1577 -1664 1627 -1647
rect 1469 -1681 1485 -1664
rect 1353 -1697 1485 -1681
rect 1611 -1681 1627 -1664
rect 1727 -1664 1777 -1647
rect 1835 -1647 2035 -1600
rect 1835 -1664 1885 -1647
rect 1727 -1681 1743 -1664
rect 1611 -1697 1743 -1681
rect 1869 -1681 1885 -1664
rect 1985 -1664 2035 -1647
rect 2093 -1647 2293 -1600
rect 2093 -1664 2143 -1647
rect 1985 -1681 2001 -1664
rect 1869 -1697 2001 -1681
rect 2127 -1681 2143 -1664
rect 2243 -1664 2293 -1647
rect 2243 -1681 2259 -1664
rect 2127 -1697 2259 -1681
<< polycont >>
rect -2243 1647 -2143 1681
rect -1985 1647 -1885 1681
rect -1727 1647 -1627 1681
rect -1469 1647 -1369 1681
rect -1211 1647 -1111 1681
rect -953 1647 -853 1681
rect -695 1647 -595 1681
rect -437 1647 -337 1681
rect -179 1647 -79 1681
rect 79 1647 179 1681
rect 337 1647 437 1681
rect 595 1647 695 1681
rect 853 1647 953 1681
rect 1111 1647 1211 1681
rect 1369 1647 1469 1681
rect 1627 1647 1727 1681
rect 1885 1647 1985 1681
rect 2143 1647 2243 1681
rect -2243 -1681 -2143 -1647
rect -1985 -1681 -1885 -1647
rect -1727 -1681 -1627 -1647
rect -1469 -1681 -1369 -1647
rect -1211 -1681 -1111 -1647
rect -953 -1681 -853 -1647
rect -695 -1681 -595 -1647
rect -437 -1681 -337 -1647
rect -179 -1681 -79 -1647
rect 79 -1681 179 -1647
rect 337 -1681 437 -1647
rect 595 -1681 695 -1647
rect 853 -1681 953 -1647
rect 1111 -1681 1211 -1647
rect 1369 -1681 1469 -1647
rect 1627 -1681 1727 -1647
rect 1885 -1681 1985 -1647
rect 2143 -1681 2243 -1647
<< locali >>
rect -2473 1785 -2377 1819
rect 2377 1785 2473 1819
rect -2473 1723 -2439 1785
rect 2439 1723 2473 1785
rect -2259 1647 -2243 1681
rect -2143 1647 -2127 1681
rect -2001 1647 -1985 1681
rect -1885 1647 -1869 1681
rect -1743 1647 -1727 1681
rect -1627 1647 -1611 1681
rect -1485 1647 -1469 1681
rect -1369 1647 -1353 1681
rect -1227 1647 -1211 1681
rect -1111 1647 -1095 1681
rect -969 1647 -953 1681
rect -853 1647 -837 1681
rect -711 1647 -695 1681
rect -595 1647 -579 1681
rect -453 1647 -437 1681
rect -337 1647 -321 1681
rect -195 1647 -179 1681
rect -79 1647 -63 1681
rect 63 1647 79 1681
rect 179 1647 195 1681
rect 321 1647 337 1681
rect 437 1647 453 1681
rect 579 1647 595 1681
rect 695 1647 711 1681
rect 837 1647 853 1681
rect 953 1647 969 1681
rect 1095 1647 1111 1681
rect 1211 1647 1227 1681
rect 1353 1647 1369 1681
rect 1469 1647 1485 1681
rect 1611 1647 1627 1681
rect 1727 1647 1743 1681
rect 1869 1647 1885 1681
rect 1985 1647 2001 1681
rect 2127 1647 2143 1681
rect 2243 1647 2259 1681
rect -2339 1588 -2305 1604
rect -2339 -1604 -2305 -1588
rect -2081 1588 -2047 1604
rect -2081 -1604 -2047 -1588
rect -1823 1588 -1789 1604
rect -1823 -1604 -1789 -1588
rect -1565 1588 -1531 1604
rect -1565 -1604 -1531 -1588
rect -1307 1588 -1273 1604
rect -1307 -1604 -1273 -1588
rect -1049 1588 -1015 1604
rect -1049 -1604 -1015 -1588
rect -791 1588 -757 1604
rect -791 -1604 -757 -1588
rect -533 1588 -499 1604
rect -533 -1604 -499 -1588
rect -275 1588 -241 1604
rect -275 -1604 -241 -1588
rect -17 1588 17 1604
rect -17 -1604 17 -1588
rect 241 1588 275 1604
rect 241 -1604 275 -1588
rect 499 1588 533 1604
rect 499 -1604 533 -1588
rect 757 1588 791 1604
rect 757 -1604 791 -1588
rect 1015 1588 1049 1604
rect 1015 -1604 1049 -1588
rect 1273 1588 1307 1604
rect 1273 -1604 1307 -1588
rect 1531 1588 1565 1604
rect 1531 -1604 1565 -1588
rect 1789 1588 1823 1604
rect 1789 -1604 1823 -1588
rect 2047 1588 2081 1604
rect 2047 -1604 2081 -1588
rect 2305 1588 2339 1604
rect 2305 -1604 2339 -1588
rect -2259 -1681 -2243 -1647
rect -2143 -1681 -2127 -1647
rect -2001 -1681 -1985 -1647
rect -1885 -1681 -1869 -1647
rect -1743 -1681 -1727 -1647
rect -1627 -1681 -1611 -1647
rect -1485 -1681 -1469 -1647
rect -1369 -1681 -1353 -1647
rect -1227 -1681 -1211 -1647
rect -1111 -1681 -1095 -1647
rect -969 -1681 -953 -1647
rect -853 -1681 -837 -1647
rect -711 -1681 -695 -1647
rect -595 -1681 -579 -1647
rect -453 -1681 -437 -1647
rect -337 -1681 -321 -1647
rect -195 -1681 -179 -1647
rect -79 -1681 -63 -1647
rect 63 -1681 79 -1647
rect 179 -1681 195 -1647
rect 321 -1681 337 -1647
rect 437 -1681 453 -1647
rect 579 -1681 595 -1647
rect 695 -1681 711 -1647
rect 837 -1681 853 -1647
rect 953 -1681 969 -1647
rect 1095 -1681 1111 -1647
rect 1211 -1681 1227 -1647
rect 1353 -1681 1369 -1647
rect 1469 -1681 1485 -1647
rect 1611 -1681 1627 -1647
rect 1727 -1681 1743 -1647
rect 1869 -1681 1885 -1647
rect 1985 -1681 2001 -1647
rect 2127 -1681 2143 -1647
rect 2243 -1681 2259 -1647
rect -2473 -1785 -2439 -1723
rect 2439 -1785 2473 -1723
rect -2473 -1819 -2377 -1785
rect 2377 -1819 2473 -1785
<< viali >>
rect -2243 1647 -2143 1681
rect -1985 1647 -1885 1681
rect -1727 1647 -1627 1681
rect -1469 1647 -1369 1681
rect -1211 1647 -1111 1681
rect -953 1647 -853 1681
rect -695 1647 -595 1681
rect -437 1647 -337 1681
rect -179 1647 -79 1681
rect 79 1647 179 1681
rect 337 1647 437 1681
rect 595 1647 695 1681
rect 853 1647 953 1681
rect 1111 1647 1211 1681
rect 1369 1647 1469 1681
rect 1627 1647 1727 1681
rect 1885 1647 1985 1681
rect 2143 1647 2243 1681
rect -2339 -1588 -2305 1588
rect -2081 -1588 -2047 1588
rect -1823 -1588 -1789 1588
rect -1565 -1588 -1531 1588
rect -1307 -1588 -1273 1588
rect -1049 -1588 -1015 1588
rect -791 -1588 -757 1588
rect -533 -1588 -499 1588
rect -275 -1588 -241 1588
rect -17 -1588 17 1588
rect 241 -1588 275 1588
rect 499 -1588 533 1588
rect 757 -1588 791 1588
rect 1015 -1588 1049 1588
rect 1273 -1588 1307 1588
rect 1531 -1588 1565 1588
rect 1789 -1588 1823 1588
rect 2047 -1588 2081 1588
rect 2305 -1588 2339 1588
rect -2243 -1681 -2143 -1647
rect -1985 -1681 -1885 -1647
rect -1727 -1681 -1627 -1647
rect -1469 -1681 -1369 -1647
rect -1211 -1681 -1111 -1647
rect -953 -1681 -853 -1647
rect -695 -1681 -595 -1647
rect -437 -1681 -337 -1647
rect -179 -1681 -79 -1647
rect 79 -1681 179 -1647
rect 337 -1681 437 -1647
rect 595 -1681 695 -1647
rect 853 -1681 953 -1647
rect 1111 -1681 1211 -1647
rect 1369 -1681 1469 -1647
rect 1627 -1681 1727 -1647
rect 1885 -1681 1985 -1647
rect 2143 -1681 2243 -1647
<< metal1 >>
rect -2255 1681 -2131 1687
rect -2255 1647 -2243 1681
rect -2143 1647 -2131 1681
rect -2255 1641 -2131 1647
rect -1997 1681 -1873 1687
rect -1997 1647 -1985 1681
rect -1885 1647 -1873 1681
rect -1997 1641 -1873 1647
rect -1739 1681 -1615 1687
rect -1739 1647 -1727 1681
rect -1627 1647 -1615 1681
rect -1739 1641 -1615 1647
rect -1481 1681 -1357 1687
rect -1481 1647 -1469 1681
rect -1369 1647 -1357 1681
rect -1481 1641 -1357 1647
rect -1223 1681 -1099 1687
rect -1223 1647 -1211 1681
rect -1111 1647 -1099 1681
rect -1223 1641 -1099 1647
rect -965 1681 -841 1687
rect -965 1647 -953 1681
rect -853 1647 -841 1681
rect -965 1641 -841 1647
rect -707 1681 -583 1687
rect -707 1647 -695 1681
rect -595 1647 -583 1681
rect -707 1641 -583 1647
rect -449 1681 -325 1687
rect -449 1647 -437 1681
rect -337 1647 -325 1681
rect -449 1641 -325 1647
rect -191 1681 -67 1687
rect -191 1647 -179 1681
rect -79 1647 -67 1681
rect -191 1641 -67 1647
rect 67 1681 191 1687
rect 67 1647 79 1681
rect 179 1647 191 1681
rect 67 1641 191 1647
rect 325 1681 449 1687
rect 325 1647 337 1681
rect 437 1647 449 1681
rect 325 1641 449 1647
rect 583 1681 707 1687
rect 583 1647 595 1681
rect 695 1647 707 1681
rect 583 1641 707 1647
rect 841 1681 965 1687
rect 841 1647 853 1681
rect 953 1647 965 1681
rect 841 1641 965 1647
rect 1099 1681 1223 1687
rect 1099 1647 1111 1681
rect 1211 1647 1223 1681
rect 1099 1641 1223 1647
rect 1357 1681 1481 1687
rect 1357 1647 1369 1681
rect 1469 1647 1481 1681
rect 1357 1641 1481 1647
rect 1615 1681 1739 1687
rect 1615 1647 1627 1681
rect 1727 1647 1739 1681
rect 1615 1641 1739 1647
rect 1873 1681 1997 1687
rect 1873 1647 1885 1681
rect 1985 1647 1997 1681
rect 1873 1641 1997 1647
rect 2131 1681 2255 1687
rect 2131 1647 2143 1681
rect 2243 1647 2255 1681
rect 2131 1641 2255 1647
rect -2345 1588 -2299 1600
rect -2345 -1588 -2339 1588
rect -2305 -1588 -2299 1588
rect -2345 -1600 -2299 -1588
rect -2087 1588 -2041 1600
rect -2087 -1588 -2081 1588
rect -2047 -1588 -2041 1588
rect -2087 -1600 -2041 -1588
rect -1829 1588 -1783 1600
rect -1829 -1588 -1823 1588
rect -1789 -1588 -1783 1588
rect -1829 -1600 -1783 -1588
rect -1571 1588 -1525 1600
rect -1571 -1588 -1565 1588
rect -1531 -1588 -1525 1588
rect -1571 -1600 -1525 -1588
rect -1313 1588 -1267 1600
rect -1313 -1588 -1307 1588
rect -1273 -1588 -1267 1588
rect -1313 -1600 -1267 -1588
rect -1055 1588 -1009 1600
rect -1055 -1588 -1049 1588
rect -1015 -1588 -1009 1588
rect -1055 -1600 -1009 -1588
rect -797 1588 -751 1600
rect -797 -1588 -791 1588
rect -757 -1588 -751 1588
rect -797 -1600 -751 -1588
rect -539 1588 -493 1600
rect -539 -1588 -533 1588
rect -499 -1588 -493 1588
rect -539 -1600 -493 -1588
rect -281 1588 -235 1600
rect -281 -1588 -275 1588
rect -241 -1588 -235 1588
rect -281 -1600 -235 -1588
rect -23 1588 23 1600
rect -23 -1588 -17 1588
rect 17 -1588 23 1588
rect -23 -1600 23 -1588
rect 235 1588 281 1600
rect 235 -1588 241 1588
rect 275 -1588 281 1588
rect 235 -1600 281 -1588
rect 493 1588 539 1600
rect 493 -1588 499 1588
rect 533 -1588 539 1588
rect 493 -1600 539 -1588
rect 751 1588 797 1600
rect 751 -1588 757 1588
rect 791 -1588 797 1588
rect 751 -1600 797 -1588
rect 1009 1588 1055 1600
rect 1009 -1588 1015 1588
rect 1049 -1588 1055 1588
rect 1009 -1600 1055 -1588
rect 1267 1588 1313 1600
rect 1267 -1588 1273 1588
rect 1307 -1588 1313 1588
rect 1267 -1600 1313 -1588
rect 1525 1588 1571 1600
rect 1525 -1588 1531 1588
rect 1565 -1588 1571 1588
rect 1525 -1600 1571 -1588
rect 1783 1588 1829 1600
rect 1783 -1588 1789 1588
rect 1823 -1588 1829 1588
rect 1783 -1600 1829 -1588
rect 2041 1588 2087 1600
rect 2041 -1588 2047 1588
rect 2081 -1588 2087 1588
rect 2041 -1600 2087 -1588
rect 2299 1588 2345 1600
rect 2299 -1588 2305 1588
rect 2339 -1588 2345 1588
rect 2299 -1600 2345 -1588
rect -2255 -1647 -2131 -1641
rect -2255 -1681 -2243 -1647
rect -2143 -1681 -2131 -1647
rect -2255 -1687 -2131 -1681
rect -1997 -1647 -1873 -1641
rect -1997 -1681 -1985 -1647
rect -1885 -1681 -1873 -1647
rect -1997 -1687 -1873 -1681
rect -1739 -1647 -1615 -1641
rect -1739 -1681 -1727 -1647
rect -1627 -1681 -1615 -1647
rect -1739 -1687 -1615 -1681
rect -1481 -1647 -1357 -1641
rect -1481 -1681 -1469 -1647
rect -1369 -1681 -1357 -1647
rect -1481 -1687 -1357 -1681
rect -1223 -1647 -1099 -1641
rect -1223 -1681 -1211 -1647
rect -1111 -1681 -1099 -1647
rect -1223 -1687 -1099 -1681
rect -965 -1647 -841 -1641
rect -965 -1681 -953 -1647
rect -853 -1681 -841 -1647
rect -965 -1687 -841 -1681
rect -707 -1647 -583 -1641
rect -707 -1681 -695 -1647
rect -595 -1681 -583 -1647
rect -707 -1687 -583 -1681
rect -449 -1647 -325 -1641
rect -449 -1681 -437 -1647
rect -337 -1681 -325 -1647
rect -449 -1687 -325 -1681
rect -191 -1647 -67 -1641
rect -191 -1681 -179 -1647
rect -79 -1681 -67 -1647
rect -191 -1687 -67 -1681
rect 67 -1647 191 -1641
rect 67 -1681 79 -1647
rect 179 -1681 191 -1647
rect 67 -1687 191 -1681
rect 325 -1647 449 -1641
rect 325 -1681 337 -1647
rect 437 -1681 449 -1647
rect 325 -1687 449 -1681
rect 583 -1647 707 -1641
rect 583 -1681 595 -1647
rect 695 -1681 707 -1647
rect 583 -1687 707 -1681
rect 841 -1647 965 -1641
rect 841 -1681 853 -1647
rect 953 -1681 965 -1647
rect 841 -1687 965 -1681
rect 1099 -1647 1223 -1641
rect 1099 -1681 1111 -1647
rect 1211 -1681 1223 -1647
rect 1099 -1687 1223 -1681
rect 1357 -1647 1481 -1641
rect 1357 -1681 1369 -1647
rect 1469 -1681 1481 -1647
rect 1357 -1687 1481 -1681
rect 1615 -1647 1739 -1641
rect 1615 -1681 1627 -1647
rect 1727 -1681 1739 -1647
rect 1615 -1687 1739 -1681
rect 1873 -1647 1997 -1641
rect 1873 -1681 1885 -1647
rect 1985 -1681 1997 -1647
rect 1873 -1687 1997 -1681
rect 2131 -1647 2255 -1641
rect 2131 -1681 2143 -1647
rect 2243 -1681 2255 -1647
rect 2131 -1687 2255 -1681
<< properties >>
string FIXED_BBOX -2456 -1802 2456 1802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 16 l 1 m 1 nf 18 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

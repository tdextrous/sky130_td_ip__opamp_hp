magic
tech sky130A
magscale 1 2
timestamp 1713234246
<< nwell >>
rect -1906 -717 1906 717
<< mvpmos >>
rect -1648 -420 -1448 420
rect -1390 -420 -1190 420
rect -1132 -420 -932 420
rect -874 -420 -674 420
rect -616 -420 -416 420
rect -358 -420 -158 420
rect -100 -420 100 420
rect 158 -420 358 420
rect 416 -420 616 420
rect 674 -420 874 420
rect 932 -420 1132 420
rect 1190 -420 1390 420
rect 1448 -420 1648 420
<< mvpdiff >>
rect -1706 408 -1648 420
rect -1706 -408 -1694 408
rect -1660 -408 -1648 408
rect -1706 -420 -1648 -408
rect -1448 408 -1390 420
rect -1448 -408 -1436 408
rect -1402 -408 -1390 408
rect -1448 -420 -1390 -408
rect -1190 408 -1132 420
rect -1190 -408 -1178 408
rect -1144 -408 -1132 408
rect -1190 -420 -1132 -408
rect -932 408 -874 420
rect -932 -408 -920 408
rect -886 -408 -874 408
rect -932 -420 -874 -408
rect -674 408 -616 420
rect -674 -408 -662 408
rect -628 -408 -616 408
rect -674 -420 -616 -408
rect -416 408 -358 420
rect -416 -408 -404 408
rect -370 -408 -358 408
rect -416 -420 -358 -408
rect -158 408 -100 420
rect -158 -408 -146 408
rect -112 -408 -100 408
rect -158 -420 -100 -408
rect 100 408 158 420
rect 100 -408 112 408
rect 146 -408 158 408
rect 100 -420 158 -408
rect 358 408 416 420
rect 358 -408 370 408
rect 404 -408 416 408
rect 358 -420 416 -408
rect 616 408 674 420
rect 616 -408 628 408
rect 662 -408 674 408
rect 616 -420 674 -408
rect 874 408 932 420
rect 874 -408 886 408
rect 920 -408 932 408
rect 874 -420 932 -408
rect 1132 408 1190 420
rect 1132 -408 1144 408
rect 1178 -408 1190 408
rect 1132 -420 1190 -408
rect 1390 408 1448 420
rect 1390 -408 1402 408
rect 1436 -408 1448 408
rect 1390 -420 1448 -408
rect 1648 408 1706 420
rect 1648 -408 1660 408
rect 1694 -408 1706 408
rect 1648 -420 1706 -408
<< mvpdiffc >>
rect -1694 -408 -1660 408
rect -1436 -408 -1402 408
rect -1178 -408 -1144 408
rect -920 -408 -886 408
rect -662 -408 -628 408
rect -404 -408 -370 408
rect -146 -408 -112 408
rect 112 -408 146 408
rect 370 -408 404 408
rect 628 -408 662 408
rect 886 -408 920 408
rect 1144 -408 1178 408
rect 1402 -408 1436 408
rect 1660 -408 1694 408
<< mvnsubdiff >>
rect -1840 639 1840 651
rect -1840 605 -1732 639
rect 1732 605 1840 639
rect -1840 593 1840 605
rect -1840 543 -1782 593
rect -1840 -543 -1828 543
rect -1794 -543 -1782 543
rect 1782 543 1840 593
rect -1840 -593 -1782 -543
rect 1782 -543 1794 543
rect 1828 -543 1840 543
rect 1782 -593 1840 -543
rect -1840 -605 1840 -593
rect -1840 -639 -1732 -605
rect 1732 -639 1840 -605
rect -1840 -651 1840 -639
<< mvnsubdiffcont >>
rect -1732 605 1732 639
rect -1828 -543 -1794 543
rect 1794 -543 1828 543
rect -1732 -639 1732 -605
<< poly >>
rect -1648 501 -1448 517
rect -1648 467 -1632 501
rect -1464 467 -1448 501
rect -1648 420 -1448 467
rect -1390 501 -1190 517
rect -1390 467 -1374 501
rect -1206 467 -1190 501
rect -1390 420 -1190 467
rect -1132 501 -932 517
rect -1132 467 -1116 501
rect -948 467 -932 501
rect -1132 420 -932 467
rect -874 501 -674 517
rect -874 467 -858 501
rect -690 467 -674 501
rect -874 420 -674 467
rect -616 501 -416 517
rect -616 467 -600 501
rect -432 467 -416 501
rect -616 420 -416 467
rect -358 501 -158 517
rect -358 467 -342 501
rect -174 467 -158 501
rect -358 420 -158 467
rect -100 501 100 517
rect -100 467 -84 501
rect 84 467 100 501
rect -100 420 100 467
rect 158 501 358 517
rect 158 467 174 501
rect 342 467 358 501
rect 158 420 358 467
rect 416 501 616 517
rect 416 467 432 501
rect 600 467 616 501
rect 416 420 616 467
rect 674 501 874 517
rect 674 467 690 501
rect 858 467 874 501
rect 674 420 874 467
rect 932 501 1132 517
rect 932 467 948 501
rect 1116 467 1132 501
rect 932 420 1132 467
rect 1190 501 1390 517
rect 1190 467 1206 501
rect 1374 467 1390 501
rect 1190 420 1390 467
rect 1448 501 1648 517
rect 1448 467 1464 501
rect 1632 467 1648 501
rect 1448 420 1648 467
rect -1648 -467 -1448 -420
rect -1648 -501 -1632 -467
rect -1464 -501 -1448 -467
rect -1648 -517 -1448 -501
rect -1390 -467 -1190 -420
rect -1390 -501 -1374 -467
rect -1206 -501 -1190 -467
rect -1390 -517 -1190 -501
rect -1132 -467 -932 -420
rect -1132 -501 -1116 -467
rect -948 -501 -932 -467
rect -1132 -517 -932 -501
rect -874 -467 -674 -420
rect -874 -501 -858 -467
rect -690 -501 -674 -467
rect -874 -517 -674 -501
rect -616 -467 -416 -420
rect -616 -501 -600 -467
rect -432 -501 -416 -467
rect -616 -517 -416 -501
rect -358 -467 -158 -420
rect -358 -501 -342 -467
rect -174 -501 -158 -467
rect -358 -517 -158 -501
rect -100 -467 100 -420
rect -100 -501 -84 -467
rect 84 -501 100 -467
rect -100 -517 100 -501
rect 158 -467 358 -420
rect 158 -501 174 -467
rect 342 -501 358 -467
rect 158 -517 358 -501
rect 416 -467 616 -420
rect 416 -501 432 -467
rect 600 -501 616 -467
rect 416 -517 616 -501
rect 674 -467 874 -420
rect 674 -501 690 -467
rect 858 -501 874 -467
rect 674 -517 874 -501
rect 932 -467 1132 -420
rect 932 -501 948 -467
rect 1116 -501 1132 -467
rect 932 -517 1132 -501
rect 1190 -467 1390 -420
rect 1190 -501 1206 -467
rect 1374 -501 1390 -467
rect 1190 -517 1390 -501
rect 1448 -467 1648 -420
rect 1448 -501 1464 -467
rect 1632 -501 1648 -467
rect 1448 -517 1648 -501
<< polycont >>
rect -1632 467 -1464 501
rect -1374 467 -1206 501
rect -1116 467 -948 501
rect -858 467 -690 501
rect -600 467 -432 501
rect -342 467 -174 501
rect -84 467 84 501
rect 174 467 342 501
rect 432 467 600 501
rect 690 467 858 501
rect 948 467 1116 501
rect 1206 467 1374 501
rect 1464 467 1632 501
rect -1632 -501 -1464 -467
rect -1374 -501 -1206 -467
rect -1116 -501 -948 -467
rect -858 -501 -690 -467
rect -600 -501 -432 -467
rect -342 -501 -174 -467
rect -84 -501 84 -467
rect 174 -501 342 -467
rect 432 -501 600 -467
rect 690 -501 858 -467
rect 948 -501 1116 -467
rect 1206 -501 1374 -467
rect 1464 -501 1632 -467
<< locali >>
rect -1828 605 -1732 639
rect 1732 605 1828 639
rect -1828 543 -1794 605
rect 1794 543 1828 605
rect -1648 467 -1632 501
rect -1464 467 -1448 501
rect -1390 467 -1374 501
rect -1206 467 -1190 501
rect -1132 467 -1116 501
rect -948 467 -932 501
rect -874 467 -858 501
rect -690 467 -674 501
rect -616 467 -600 501
rect -432 467 -416 501
rect -358 467 -342 501
rect -174 467 -158 501
rect -100 467 -84 501
rect 84 467 100 501
rect 158 467 174 501
rect 342 467 358 501
rect 416 467 432 501
rect 600 467 616 501
rect 674 467 690 501
rect 858 467 874 501
rect 932 467 948 501
rect 1116 467 1132 501
rect 1190 467 1206 501
rect 1374 467 1390 501
rect 1448 467 1464 501
rect 1632 467 1648 501
rect -1694 408 -1660 424
rect -1694 -424 -1660 -408
rect -1436 408 -1402 424
rect -1436 -424 -1402 -408
rect -1178 408 -1144 424
rect -1178 -424 -1144 -408
rect -920 408 -886 424
rect -920 -424 -886 -408
rect -662 408 -628 424
rect -662 -424 -628 -408
rect -404 408 -370 424
rect -404 -424 -370 -408
rect -146 408 -112 424
rect -146 -424 -112 -408
rect 112 408 146 424
rect 112 -424 146 -408
rect 370 408 404 424
rect 370 -424 404 -408
rect 628 408 662 424
rect 628 -424 662 -408
rect 886 408 920 424
rect 886 -424 920 -408
rect 1144 408 1178 424
rect 1144 -424 1178 -408
rect 1402 408 1436 424
rect 1402 -424 1436 -408
rect 1660 408 1694 424
rect 1660 -424 1694 -408
rect -1648 -501 -1632 -467
rect -1464 -501 -1448 -467
rect -1390 -501 -1374 -467
rect -1206 -501 -1190 -467
rect -1132 -501 -1116 -467
rect -948 -501 -932 -467
rect -874 -501 -858 -467
rect -690 -501 -674 -467
rect -616 -501 -600 -467
rect -432 -501 -416 -467
rect -358 -501 -342 -467
rect -174 -501 -158 -467
rect -100 -501 -84 -467
rect 84 -501 100 -467
rect 158 -501 174 -467
rect 342 -501 358 -467
rect 416 -501 432 -467
rect 600 -501 616 -467
rect 674 -501 690 -467
rect 858 -501 874 -467
rect 932 -501 948 -467
rect 1116 -501 1132 -467
rect 1190 -501 1206 -467
rect 1374 -501 1390 -467
rect 1448 -501 1464 -467
rect 1632 -501 1648 -467
rect -1828 -605 -1794 -543
rect 1794 -605 1828 -543
rect -1828 -639 -1732 -605
rect 1732 -639 1828 -605
<< viali >>
rect -1632 467 -1464 501
rect -1374 467 -1206 501
rect -1116 467 -948 501
rect -858 467 -690 501
rect -600 467 -432 501
rect -342 467 -174 501
rect -84 467 84 501
rect 174 467 342 501
rect 432 467 600 501
rect 690 467 858 501
rect 948 467 1116 501
rect 1206 467 1374 501
rect 1464 467 1632 501
rect -1694 -408 -1660 408
rect -1436 -408 -1402 408
rect -1178 -408 -1144 408
rect -920 -408 -886 408
rect -662 -408 -628 408
rect -404 -408 -370 408
rect -146 -408 -112 408
rect 112 -408 146 408
rect 370 -408 404 408
rect 628 -408 662 408
rect 886 -408 920 408
rect 1144 -408 1178 408
rect 1402 -408 1436 408
rect 1660 -408 1694 408
rect -1632 -501 -1464 -467
rect -1374 -501 -1206 -467
rect -1116 -501 -948 -467
rect -858 -501 -690 -467
rect -600 -501 -432 -467
rect -342 -501 -174 -467
rect -84 -501 84 -467
rect 174 -501 342 -467
rect 432 -501 600 -467
rect 690 -501 858 -467
rect 948 -501 1116 -467
rect 1206 -501 1374 -467
rect 1464 -501 1632 -467
<< metal1 >>
rect -1644 501 -1452 507
rect -1644 467 -1632 501
rect -1464 467 -1452 501
rect -1644 461 -1452 467
rect -1386 501 -1194 507
rect -1386 467 -1374 501
rect -1206 467 -1194 501
rect -1386 461 -1194 467
rect -1128 501 -936 507
rect -1128 467 -1116 501
rect -948 467 -936 501
rect -1128 461 -936 467
rect -870 501 -678 507
rect -870 467 -858 501
rect -690 467 -678 501
rect -870 461 -678 467
rect -612 501 -420 507
rect -612 467 -600 501
rect -432 467 -420 501
rect -612 461 -420 467
rect -354 501 -162 507
rect -354 467 -342 501
rect -174 467 -162 501
rect -354 461 -162 467
rect -96 501 96 507
rect -96 467 -84 501
rect 84 467 96 501
rect -96 461 96 467
rect 162 501 354 507
rect 162 467 174 501
rect 342 467 354 501
rect 162 461 354 467
rect 420 501 612 507
rect 420 467 432 501
rect 600 467 612 501
rect 420 461 612 467
rect 678 501 870 507
rect 678 467 690 501
rect 858 467 870 501
rect 678 461 870 467
rect 936 501 1128 507
rect 936 467 948 501
rect 1116 467 1128 501
rect 936 461 1128 467
rect 1194 501 1386 507
rect 1194 467 1206 501
rect 1374 467 1386 501
rect 1194 461 1386 467
rect 1452 501 1644 507
rect 1452 467 1464 501
rect 1632 467 1644 501
rect 1452 461 1644 467
rect -1700 408 -1654 420
rect -1700 -408 -1694 408
rect -1660 -408 -1654 408
rect -1700 -420 -1654 -408
rect -1442 408 -1396 420
rect -1442 -408 -1436 408
rect -1402 -408 -1396 408
rect -1442 -420 -1396 -408
rect -1184 408 -1138 420
rect -1184 -408 -1178 408
rect -1144 -408 -1138 408
rect -1184 -420 -1138 -408
rect -926 408 -880 420
rect -926 -408 -920 408
rect -886 -408 -880 408
rect -926 -420 -880 -408
rect -668 408 -622 420
rect -668 -408 -662 408
rect -628 -408 -622 408
rect -668 -420 -622 -408
rect -410 408 -364 420
rect -410 -408 -404 408
rect -370 -408 -364 408
rect -410 -420 -364 -408
rect -152 408 -106 420
rect -152 -408 -146 408
rect -112 -408 -106 408
rect -152 -420 -106 -408
rect 106 408 152 420
rect 106 -408 112 408
rect 146 -408 152 408
rect 106 -420 152 -408
rect 364 408 410 420
rect 364 -408 370 408
rect 404 -408 410 408
rect 364 -420 410 -408
rect 622 408 668 420
rect 622 -408 628 408
rect 662 -408 668 408
rect 622 -420 668 -408
rect 880 408 926 420
rect 880 -408 886 408
rect 920 -408 926 408
rect 880 -420 926 -408
rect 1138 408 1184 420
rect 1138 -408 1144 408
rect 1178 -408 1184 408
rect 1138 -420 1184 -408
rect 1396 408 1442 420
rect 1396 -408 1402 408
rect 1436 -408 1442 408
rect 1396 -420 1442 -408
rect 1654 408 1700 420
rect 1654 -408 1660 408
rect 1694 -408 1700 408
rect 1654 -420 1700 -408
rect -1644 -467 -1452 -461
rect -1644 -501 -1632 -467
rect -1464 -501 -1452 -467
rect -1644 -507 -1452 -501
rect -1386 -467 -1194 -461
rect -1386 -501 -1374 -467
rect -1206 -501 -1194 -467
rect -1386 -507 -1194 -501
rect -1128 -467 -936 -461
rect -1128 -501 -1116 -467
rect -948 -501 -936 -467
rect -1128 -507 -936 -501
rect -870 -467 -678 -461
rect -870 -501 -858 -467
rect -690 -501 -678 -467
rect -870 -507 -678 -501
rect -612 -467 -420 -461
rect -612 -501 -600 -467
rect -432 -501 -420 -467
rect -612 -507 -420 -501
rect -354 -467 -162 -461
rect -354 -501 -342 -467
rect -174 -501 -162 -467
rect -354 -507 -162 -501
rect -96 -467 96 -461
rect -96 -501 -84 -467
rect 84 -501 96 -467
rect -96 -507 96 -501
rect 162 -467 354 -461
rect 162 -501 174 -467
rect 342 -501 354 -467
rect 162 -507 354 -501
rect 420 -467 612 -461
rect 420 -501 432 -467
rect 600 -501 612 -467
rect 420 -507 612 -501
rect 678 -467 870 -461
rect 678 -501 690 -467
rect 858 -501 870 -467
rect 678 -507 870 -501
rect 936 -467 1128 -461
rect 936 -501 948 -467
rect 1116 -501 1128 -467
rect 936 -507 1128 -501
rect 1194 -467 1386 -461
rect 1194 -501 1206 -467
rect 1374 -501 1386 -467
rect 1194 -507 1386 -501
rect 1452 -467 1644 -461
rect 1452 -501 1464 -467
rect 1632 -501 1644 -467
rect 1452 -507 1644 -501
<< properties >>
string FIXED_BBOX -1811 -622 1811 622
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.2 l 1 m 1 nf 13 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713234246
<< nwell >>
rect -4615 -2797 4615 2797
<< mvpmos >>
rect -4357 -2500 -4157 2500
rect -4099 -2500 -3899 2500
rect -3841 -2500 -3641 2500
rect -3583 -2500 -3383 2500
rect -3325 -2500 -3125 2500
rect -3067 -2500 -2867 2500
rect -2809 -2500 -2609 2500
rect -2551 -2500 -2351 2500
rect -2293 -2500 -2093 2500
rect -2035 -2500 -1835 2500
rect -1777 -2500 -1577 2500
rect -1519 -2500 -1319 2500
rect -1261 -2500 -1061 2500
rect -1003 -2500 -803 2500
rect -745 -2500 -545 2500
rect -487 -2500 -287 2500
rect -229 -2500 -29 2500
rect 29 -2500 229 2500
rect 287 -2500 487 2500
rect 545 -2500 745 2500
rect 803 -2500 1003 2500
rect 1061 -2500 1261 2500
rect 1319 -2500 1519 2500
rect 1577 -2500 1777 2500
rect 1835 -2500 2035 2500
rect 2093 -2500 2293 2500
rect 2351 -2500 2551 2500
rect 2609 -2500 2809 2500
rect 2867 -2500 3067 2500
rect 3125 -2500 3325 2500
rect 3383 -2500 3583 2500
rect 3641 -2500 3841 2500
rect 3899 -2500 4099 2500
rect 4157 -2500 4357 2500
<< mvpdiff >>
rect -4415 2488 -4357 2500
rect -4415 -2488 -4403 2488
rect -4369 -2488 -4357 2488
rect -4415 -2500 -4357 -2488
rect -4157 2488 -4099 2500
rect -4157 -2488 -4145 2488
rect -4111 -2488 -4099 2488
rect -4157 -2500 -4099 -2488
rect -3899 2488 -3841 2500
rect -3899 -2488 -3887 2488
rect -3853 -2488 -3841 2488
rect -3899 -2500 -3841 -2488
rect -3641 2488 -3583 2500
rect -3641 -2488 -3629 2488
rect -3595 -2488 -3583 2488
rect -3641 -2500 -3583 -2488
rect -3383 2488 -3325 2500
rect -3383 -2488 -3371 2488
rect -3337 -2488 -3325 2488
rect -3383 -2500 -3325 -2488
rect -3125 2488 -3067 2500
rect -3125 -2488 -3113 2488
rect -3079 -2488 -3067 2488
rect -3125 -2500 -3067 -2488
rect -2867 2488 -2809 2500
rect -2867 -2488 -2855 2488
rect -2821 -2488 -2809 2488
rect -2867 -2500 -2809 -2488
rect -2609 2488 -2551 2500
rect -2609 -2488 -2597 2488
rect -2563 -2488 -2551 2488
rect -2609 -2500 -2551 -2488
rect -2351 2488 -2293 2500
rect -2351 -2488 -2339 2488
rect -2305 -2488 -2293 2488
rect -2351 -2500 -2293 -2488
rect -2093 2488 -2035 2500
rect -2093 -2488 -2081 2488
rect -2047 -2488 -2035 2488
rect -2093 -2500 -2035 -2488
rect -1835 2488 -1777 2500
rect -1835 -2488 -1823 2488
rect -1789 -2488 -1777 2488
rect -1835 -2500 -1777 -2488
rect -1577 2488 -1519 2500
rect -1577 -2488 -1565 2488
rect -1531 -2488 -1519 2488
rect -1577 -2500 -1519 -2488
rect -1319 2488 -1261 2500
rect -1319 -2488 -1307 2488
rect -1273 -2488 -1261 2488
rect -1319 -2500 -1261 -2488
rect -1061 2488 -1003 2500
rect -1061 -2488 -1049 2488
rect -1015 -2488 -1003 2488
rect -1061 -2500 -1003 -2488
rect -803 2488 -745 2500
rect -803 -2488 -791 2488
rect -757 -2488 -745 2488
rect -803 -2500 -745 -2488
rect -545 2488 -487 2500
rect -545 -2488 -533 2488
rect -499 -2488 -487 2488
rect -545 -2500 -487 -2488
rect -287 2488 -229 2500
rect -287 -2488 -275 2488
rect -241 -2488 -229 2488
rect -287 -2500 -229 -2488
rect -29 2488 29 2500
rect -29 -2488 -17 2488
rect 17 -2488 29 2488
rect -29 -2500 29 -2488
rect 229 2488 287 2500
rect 229 -2488 241 2488
rect 275 -2488 287 2488
rect 229 -2500 287 -2488
rect 487 2488 545 2500
rect 487 -2488 499 2488
rect 533 -2488 545 2488
rect 487 -2500 545 -2488
rect 745 2488 803 2500
rect 745 -2488 757 2488
rect 791 -2488 803 2488
rect 745 -2500 803 -2488
rect 1003 2488 1061 2500
rect 1003 -2488 1015 2488
rect 1049 -2488 1061 2488
rect 1003 -2500 1061 -2488
rect 1261 2488 1319 2500
rect 1261 -2488 1273 2488
rect 1307 -2488 1319 2488
rect 1261 -2500 1319 -2488
rect 1519 2488 1577 2500
rect 1519 -2488 1531 2488
rect 1565 -2488 1577 2488
rect 1519 -2500 1577 -2488
rect 1777 2488 1835 2500
rect 1777 -2488 1789 2488
rect 1823 -2488 1835 2488
rect 1777 -2500 1835 -2488
rect 2035 2488 2093 2500
rect 2035 -2488 2047 2488
rect 2081 -2488 2093 2488
rect 2035 -2500 2093 -2488
rect 2293 2488 2351 2500
rect 2293 -2488 2305 2488
rect 2339 -2488 2351 2488
rect 2293 -2500 2351 -2488
rect 2551 2488 2609 2500
rect 2551 -2488 2563 2488
rect 2597 -2488 2609 2488
rect 2551 -2500 2609 -2488
rect 2809 2488 2867 2500
rect 2809 -2488 2821 2488
rect 2855 -2488 2867 2488
rect 2809 -2500 2867 -2488
rect 3067 2488 3125 2500
rect 3067 -2488 3079 2488
rect 3113 -2488 3125 2488
rect 3067 -2500 3125 -2488
rect 3325 2488 3383 2500
rect 3325 -2488 3337 2488
rect 3371 -2488 3383 2488
rect 3325 -2500 3383 -2488
rect 3583 2488 3641 2500
rect 3583 -2488 3595 2488
rect 3629 -2488 3641 2488
rect 3583 -2500 3641 -2488
rect 3841 2488 3899 2500
rect 3841 -2488 3853 2488
rect 3887 -2488 3899 2488
rect 3841 -2500 3899 -2488
rect 4099 2488 4157 2500
rect 4099 -2488 4111 2488
rect 4145 -2488 4157 2488
rect 4099 -2500 4157 -2488
rect 4357 2488 4415 2500
rect 4357 -2488 4369 2488
rect 4403 -2488 4415 2488
rect 4357 -2500 4415 -2488
<< mvpdiffc >>
rect -4403 -2488 -4369 2488
rect -4145 -2488 -4111 2488
rect -3887 -2488 -3853 2488
rect -3629 -2488 -3595 2488
rect -3371 -2488 -3337 2488
rect -3113 -2488 -3079 2488
rect -2855 -2488 -2821 2488
rect -2597 -2488 -2563 2488
rect -2339 -2488 -2305 2488
rect -2081 -2488 -2047 2488
rect -1823 -2488 -1789 2488
rect -1565 -2488 -1531 2488
rect -1307 -2488 -1273 2488
rect -1049 -2488 -1015 2488
rect -791 -2488 -757 2488
rect -533 -2488 -499 2488
rect -275 -2488 -241 2488
rect -17 -2488 17 2488
rect 241 -2488 275 2488
rect 499 -2488 533 2488
rect 757 -2488 791 2488
rect 1015 -2488 1049 2488
rect 1273 -2488 1307 2488
rect 1531 -2488 1565 2488
rect 1789 -2488 1823 2488
rect 2047 -2488 2081 2488
rect 2305 -2488 2339 2488
rect 2563 -2488 2597 2488
rect 2821 -2488 2855 2488
rect 3079 -2488 3113 2488
rect 3337 -2488 3371 2488
rect 3595 -2488 3629 2488
rect 3853 -2488 3887 2488
rect 4111 -2488 4145 2488
rect 4369 -2488 4403 2488
<< mvnsubdiff >>
rect -4549 2719 4549 2731
rect -4549 2685 -4441 2719
rect 4441 2685 4549 2719
rect -4549 2673 4549 2685
rect -4549 2623 -4491 2673
rect -4549 -2623 -4537 2623
rect -4503 -2623 -4491 2623
rect 4491 2623 4549 2673
rect -4549 -2673 -4491 -2623
rect 4491 -2623 4503 2623
rect 4537 -2623 4549 2623
rect 4491 -2673 4549 -2623
rect -4549 -2685 4549 -2673
rect -4549 -2719 -4441 -2685
rect 4441 -2719 4549 -2685
rect -4549 -2731 4549 -2719
<< mvnsubdiffcont >>
rect -4441 2685 4441 2719
rect -4537 -2623 -4503 2623
rect 4503 -2623 4537 2623
rect -4441 -2719 4441 -2685
<< poly >>
rect -4357 2581 -4157 2597
rect -4357 2547 -4341 2581
rect -4173 2547 -4157 2581
rect -4357 2500 -4157 2547
rect -4099 2581 -3899 2597
rect -4099 2547 -4083 2581
rect -3915 2547 -3899 2581
rect -4099 2500 -3899 2547
rect -3841 2581 -3641 2597
rect -3841 2547 -3825 2581
rect -3657 2547 -3641 2581
rect -3841 2500 -3641 2547
rect -3583 2581 -3383 2597
rect -3583 2547 -3567 2581
rect -3399 2547 -3383 2581
rect -3583 2500 -3383 2547
rect -3325 2581 -3125 2597
rect -3325 2547 -3309 2581
rect -3141 2547 -3125 2581
rect -3325 2500 -3125 2547
rect -3067 2581 -2867 2597
rect -3067 2547 -3051 2581
rect -2883 2547 -2867 2581
rect -3067 2500 -2867 2547
rect -2809 2581 -2609 2597
rect -2809 2547 -2793 2581
rect -2625 2547 -2609 2581
rect -2809 2500 -2609 2547
rect -2551 2581 -2351 2597
rect -2551 2547 -2535 2581
rect -2367 2547 -2351 2581
rect -2551 2500 -2351 2547
rect -2293 2581 -2093 2597
rect -2293 2547 -2277 2581
rect -2109 2547 -2093 2581
rect -2293 2500 -2093 2547
rect -2035 2581 -1835 2597
rect -2035 2547 -2019 2581
rect -1851 2547 -1835 2581
rect -2035 2500 -1835 2547
rect -1777 2581 -1577 2597
rect -1777 2547 -1761 2581
rect -1593 2547 -1577 2581
rect -1777 2500 -1577 2547
rect -1519 2581 -1319 2597
rect -1519 2547 -1503 2581
rect -1335 2547 -1319 2581
rect -1519 2500 -1319 2547
rect -1261 2581 -1061 2597
rect -1261 2547 -1245 2581
rect -1077 2547 -1061 2581
rect -1261 2500 -1061 2547
rect -1003 2581 -803 2597
rect -1003 2547 -987 2581
rect -819 2547 -803 2581
rect -1003 2500 -803 2547
rect -745 2581 -545 2597
rect -745 2547 -729 2581
rect -561 2547 -545 2581
rect -745 2500 -545 2547
rect -487 2581 -287 2597
rect -487 2547 -471 2581
rect -303 2547 -287 2581
rect -487 2500 -287 2547
rect -229 2581 -29 2597
rect -229 2547 -213 2581
rect -45 2547 -29 2581
rect -229 2500 -29 2547
rect 29 2581 229 2597
rect 29 2547 45 2581
rect 213 2547 229 2581
rect 29 2500 229 2547
rect 287 2581 487 2597
rect 287 2547 303 2581
rect 471 2547 487 2581
rect 287 2500 487 2547
rect 545 2581 745 2597
rect 545 2547 561 2581
rect 729 2547 745 2581
rect 545 2500 745 2547
rect 803 2581 1003 2597
rect 803 2547 819 2581
rect 987 2547 1003 2581
rect 803 2500 1003 2547
rect 1061 2581 1261 2597
rect 1061 2547 1077 2581
rect 1245 2547 1261 2581
rect 1061 2500 1261 2547
rect 1319 2581 1519 2597
rect 1319 2547 1335 2581
rect 1503 2547 1519 2581
rect 1319 2500 1519 2547
rect 1577 2581 1777 2597
rect 1577 2547 1593 2581
rect 1761 2547 1777 2581
rect 1577 2500 1777 2547
rect 1835 2581 2035 2597
rect 1835 2547 1851 2581
rect 2019 2547 2035 2581
rect 1835 2500 2035 2547
rect 2093 2581 2293 2597
rect 2093 2547 2109 2581
rect 2277 2547 2293 2581
rect 2093 2500 2293 2547
rect 2351 2581 2551 2597
rect 2351 2547 2367 2581
rect 2535 2547 2551 2581
rect 2351 2500 2551 2547
rect 2609 2581 2809 2597
rect 2609 2547 2625 2581
rect 2793 2547 2809 2581
rect 2609 2500 2809 2547
rect 2867 2581 3067 2597
rect 2867 2547 2883 2581
rect 3051 2547 3067 2581
rect 2867 2500 3067 2547
rect 3125 2581 3325 2597
rect 3125 2547 3141 2581
rect 3309 2547 3325 2581
rect 3125 2500 3325 2547
rect 3383 2581 3583 2597
rect 3383 2547 3399 2581
rect 3567 2547 3583 2581
rect 3383 2500 3583 2547
rect 3641 2581 3841 2597
rect 3641 2547 3657 2581
rect 3825 2547 3841 2581
rect 3641 2500 3841 2547
rect 3899 2581 4099 2597
rect 3899 2547 3915 2581
rect 4083 2547 4099 2581
rect 3899 2500 4099 2547
rect 4157 2581 4357 2597
rect 4157 2547 4173 2581
rect 4341 2547 4357 2581
rect 4157 2500 4357 2547
rect -4357 -2547 -4157 -2500
rect -4357 -2581 -4341 -2547
rect -4173 -2581 -4157 -2547
rect -4357 -2597 -4157 -2581
rect -4099 -2547 -3899 -2500
rect -4099 -2581 -4083 -2547
rect -3915 -2581 -3899 -2547
rect -4099 -2597 -3899 -2581
rect -3841 -2547 -3641 -2500
rect -3841 -2581 -3825 -2547
rect -3657 -2581 -3641 -2547
rect -3841 -2597 -3641 -2581
rect -3583 -2547 -3383 -2500
rect -3583 -2581 -3567 -2547
rect -3399 -2581 -3383 -2547
rect -3583 -2597 -3383 -2581
rect -3325 -2547 -3125 -2500
rect -3325 -2581 -3309 -2547
rect -3141 -2581 -3125 -2547
rect -3325 -2597 -3125 -2581
rect -3067 -2547 -2867 -2500
rect -3067 -2581 -3051 -2547
rect -2883 -2581 -2867 -2547
rect -3067 -2597 -2867 -2581
rect -2809 -2547 -2609 -2500
rect -2809 -2581 -2793 -2547
rect -2625 -2581 -2609 -2547
rect -2809 -2597 -2609 -2581
rect -2551 -2547 -2351 -2500
rect -2551 -2581 -2535 -2547
rect -2367 -2581 -2351 -2547
rect -2551 -2597 -2351 -2581
rect -2293 -2547 -2093 -2500
rect -2293 -2581 -2277 -2547
rect -2109 -2581 -2093 -2547
rect -2293 -2597 -2093 -2581
rect -2035 -2547 -1835 -2500
rect -2035 -2581 -2019 -2547
rect -1851 -2581 -1835 -2547
rect -2035 -2597 -1835 -2581
rect -1777 -2547 -1577 -2500
rect -1777 -2581 -1761 -2547
rect -1593 -2581 -1577 -2547
rect -1777 -2597 -1577 -2581
rect -1519 -2547 -1319 -2500
rect -1519 -2581 -1503 -2547
rect -1335 -2581 -1319 -2547
rect -1519 -2597 -1319 -2581
rect -1261 -2547 -1061 -2500
rect -1261 -2581 -1245 -2547
rect -1077 -2581 -1061 -2547
rect -1261 -2597 -1061 -2581
rect -1003 -2547 -803 -2500
rect -1003 -2581 -987 -2547
rect -819 -2581 -803 -2547
rect -1003 -2597 -803 -2581
rect -745 -2547 -545 -2500
rect -745 -2581 -729 -2547
rect -561 -2581 -545 -2547
rect -745 -2597 -545 -2581
rect -487 -2547 -287 -2500
rect -487 -2581 -471 -2547
rect -303 -2581 -287 -2547
rect -487 -2597 -287 -2581
rect -229 -2547 -29 -2500
rect -229 -2581 -213 -2547
rect -45 -2581 -29 -2547
rect -229 -2597 -29 -2581
rect 29 -2547 229 -2500
rect 29 -2581 45 -2547
rect 213 -2581 229 -2547
rect 29 -2597 229 -2581
rect 287 -2547 487 -2500
rect 287 -2581 303 -2547
rect 471 -2581 487 -2547
rect 287 -2597 487 -2581
rect 545 -2547 745 -2500
rect 545 -2581 561 -2547
rect 729 -2581 745 -2547
rect 545 -2597 745 -2581
rect 803 -2547 1003 -2500
rect 803 -2581 819 -2547
rect 987 -2581 1003 -2547
rect 803 -2597 1003 -2581
rect 1061 -2547 1261 -2500
rect 1061 -2581 1077 -2547
rect 1245 -2581 1261 -2547
rect 1061 -2597 1261 -2581
rect 1319 -2547 1519 -2500
rect 1319 -2581 1335 -2547
rect 1503 -2581 1519 -2547
rect 1319 -2597 1519 -2581
rect 1577 -2547 1777 -2500
rect 1577 -2581 1593 -2547
rect 1761 -2581 1777 -2547
rect 1577 -2597 1777 -2581
rect 1835 -2547 2035 -2500
rect 1835 -2581 1851 -2547
rect 2019 -2581 2035 -2547
rect 1835 -2597 2035 -2581
rect 2093 -2547 2293 -2500
rect 2093 -2581 2109 -2547
rect 2277 -2581 2293 -2547
rect 2093 -2597 2293 -2581
rect 2351 -2547 2551 -2500
rect 2351 -2581 2367 -2547
rect 2535 -2581 2551 -2547
rect 2351 -2597 2551 -2581
rect 2609 -2547 2809 -2500
rect 2609 -2581 2625 -2547
rect 2793 -2581 2809 -2547
rect 2609 -2597 2809 -2581
rect 2867 -2547 3067 -2500
rect 2867 -2581 2883 -2547
rect 3051 -2581 3067 -2547
rect 2867 -2597 3067 -2581
rect 3125 -2547 3325 -2500
rect 3125 -2581 3141 -2547
rect 3309 -2581 3325 -2547
rect 3125 -2597 3325 -2581
rect 3383 -2547 3583 -2500
rect 3383 -2581 3399 -2547
rect 3567 -2581 3583 -2547
rect 3383 -2597 3583 -2581
rect 3641 -2547 3841 -2500
rect 3641 -2581 3657 -2547
rect 3825 -2581 3841 -2547
rect 3641 -2597 3841 -2581
rect 3899 -2547 4099 -2500
rect 3899 -2581 3915 -2547
rect 4083 -2581 4099 -2547
rect 3899 -2597 4099 -2581
rect 4157 -2547 4357 -2500
rect 4157 -2581 4173 -2547
rect 4341 -2581 4357 -2547
rect 4157 -2597 4357 -2581
<< polycont >>
rect -4341 2547 -4173 2581
rect -4083 2547 -3915 2581
rect -3825 2547 -3657 2581
rect -3567 2547 -3399 2581
rect -3309 2547 -3141 2581
rect -3051 2547 -2883 2581
rect -2793 2547 -2625 2581
rect -2535 2547 -2367 2581
rect -2277 2547 -2109 2581
rect -2019 2547 -1851 2581
rect -1761 2547 -1593 2581
rect -1503 2547 -1335 2581
rect -1245 2547 -1077 2581
rect -987 2547 -819 2581
rect -729 2547 -561 2581
rect -471 2547 -303 2581
rect -213 2547 -45 2581
rect 45 2547 213 2581
rect 303 2547 471 2581
rect 561 2547 729 2581
rect 819 2547 987 2581
rect 1077 2547 1245 2581
rect 1335 2547 1503 2581
rect 1593 2547 1761 2581
rect 1851 2547 2019 2581
rect 2109 2547 2277 2581
rect 2367 2547 2535 2581
rect 2625 2547 2793 2581
rect 2883 2547 3051 2581
rect 3141 2547 3309 2581
rect 3399 2547 3567 2581
rect 3657 2547 3825 2581
rect 3915 2547 4083 2581
rect 4173 2547 4341 2581
rect -4341 -2581 -4173 -2547
rect -4083 -2581 -3915 -2547
rect -3825 -2581 -3657 -2547
rect -3567 -2581 -3399 -2547
rect -3309 -2581 -3141 -2547
rect -3051 -2581 -2883 -2547
rect -2793 -2581 -2625 -2547
rect -2535 -2581 -2367 -2547
rect -2277 -2581 -2109 -2547
rect -2019 -2581 -1851 -2547
rect -1761 -2581 -1593 -2547
rect -1503 -2581 -1335 -2547
rect -1245 -2581 -1077 -2547
rect -987 -2581 -819 -2547
rect -729 -2581 -561 -2547
rect -471 -2581 -303 -2547
rect -213 -2581 -45 -2547
rect 45 -2581 213 -2547
rect 303 -2581 471 -2547
rect 561 -2581 729 -2547
rect 819 -2581 987 -2547
rect 1077 -2581 1245 -2547
rect 1335 -2581 1503 -2547
rect 1593 -2581 1761 -2547
rect 1851 -2581 2019 -2547
rect 2109 -2581 2277 -2547
rect 2367 -2581 2535 -2547
rect 2625 -2581 2793 -2547
rect 2883 -2581 3051 -2547
rect 3141 -2581 3309 -2547
rect 3399 -2581 3567 -2547
rect 3657 -2581 3825 -2547
rect 3915 -2581 4083 -2547
rect 4173 -2581 4341 -2547
<< locali >>
rect -4537 2685 -4441 2719
rect 4441 2685 4537 2719
rect -4537 2623 -4503 2685
rect 4503 2623 4537 2685
rect -4357 2547 -4341 2581
rect -4173 2547 -4157 2581
rect -4099 2547 -4083 2581
rect -3915 2547 -3899 2581
rect -3841 2547 -3825 2581
rect -3657 2547 -3641 2581
rect -3583 2547 -3567 2581
rect -3399 2547 -3383 2581
rect -3325 2547 -3309 2581
rect -3141 2547 -3125 2581
rect -3067 2547 -3051 2581
rect -2883 2547 -2867 2581
rect -2809 2547 -2793 2581
rect -2625 2547 -2609 2581
rect -2551 2547 -2535 2581
rect -2367 2547 -2351 2581
rect -2293 2547 -2277 2581
rect -2109 2547 -2093 2581
rect -2035 2547 -2019 2581
rect -1851 2547 -1835 2581
rect -1777 2547 -1761 2581
rect -1593 2547 -1577 2581
rect -1519 2547 -1503 2581
rect -1335 2547 -1319 2581
rect -1261 2547 -1245 2581
rect -1077 2547 -1061 2581
rect -1003 2547 -987 2581
rect -819 2547 -803 2581
rect -745 2547 -729 2581
rect -561 2547 -545 2581
rect -487 2547 -471 2581
rect -303 2547 -287 2581
rect -229 2547 -213 2581
rect -45 2547 -29 2581
rect 29 2547 45 2581
rect 213 2547 229 2581
rect 287 2547 303 2581
rect 471 2547 487 2581
rect 545 2547 561 2581
rect 729 2547 745 2581
rect 803 2547 819 2581
rect 987 2547 1003 2581
rect 1061 2547 1077 2581
rect 1245 2547 1261 2581
rect 1319 2547 1335 2581
rect 1503 2547 1519 2581
rect 1577 2547 1593 2581
rect 1761 2547 1777 2581
rect 1835 2547 1851 2581
rect 2019 2547 2035 2581
rect 2093 2547 2109 2581
rect 2277 2547 2293 2581
rect 2351 2547 2367 2581
rect 2535 2547 2551 2581
rect 2609 2547 2625 2581
rect 2793 2547 2809 2581
rect 2867 2547 2883 2581
rect 3051 2547 3067 2581
rect 3125 2547 3141 2581
rect 3309 2547 3325 2581
rect 3383 2547 3399 2581
rect 3567 2547 3583 2581
rect 3641 2547 3657 2581
rect 3825 2547 3841 2581
rect 3899 2547 3915 2581
rect 4083 2547 4099 2581
rect 4157 2547 4173 2581
rect 4341 2547 4357 2581
rect -4403 2488 -4369 2504
rect -4403 -2504 -4369 -2488
rect -4145 2488 -4111 2504
rect -4145 -2504 -4111 -2488
rect -3887 2488 -3853 2504
rect -3887 -2504 -3853 -2488
rect -3629 2488 -3595 2504
rect -3629 -2504 -3595 -2488
rect -3371 2488 -3337 2504
rect -3371 -2504 -3337 -2488
rect -3113 2488 -3079 2504
rect -3113 -2504 -3079 -2488
rect -2855 2488 -2821 2504
rect -2855 -2504 -2821 -2488
rect -2597 2488 -2563 2504
rect -2597 -2504 -2563 -2488
rect -2339 2488 -2305 2504
rect -2339 -2504 -2305 -2488
rect -2081 2488 -2047 2504
rect -2081 -2504 -2047 -2488
rect -1823 2488 -1789 2504
rect -1823 -2504 -1789 -2488
rect -1565 2488 -1531 2504
rect -1565 -2504 -1531 -2488
rect -1307 2488 -1273 2504
rect -1307 -2504 -1273 -2488
rect -1049 2488 -1015 2504
rect -1049 -2504 -1015 -2488
rect -791 2488 -757 2504
rect -791 -2504 -757 -2488
rect -533 2488 -499 2504
rect -533 -2504 -499 -2488
rect -275 2488 -241 2504
rect -275 -2504 -241 -2488
rect -17 2488 17 2504
rect -17 -2504 17 -2488
rect 241 2488 275 2504
rect 241 -2504 275 -2488
rect 499 2488 533 2504
rect 499 -2504 533 -2488
rect 757 2488 791 2504
rect 757 -2504 791 -2488
rect 1015 2488 1049 2504
rect 1015 -2504 1049 -2488
rect 1273 2488 1307 2504
rect 1273 -2504 1307 -2488
rect 1531 2488 1565 2504
rect 1531 -2504 1565 -2488
rect 1789 2488 1823 2504
rect 1789 -2504 1823 -2488
rect 2047 2488 2081 2504
rect 2047 -2504 2081 -2488
rect 2305 2488 2339 2504
rect 2305 -2504 2339 -2488
rect 2563 2488 2597 2504
rect 2563 -2504 2597 -2488
rect 2821 2488 2855 2504
rect 2821 -2504 2855 -2488
rect 3079 2488 3113 2504
rect 3079 -2504 3113 -2488
rect 3337 2488 3371 2504
rect 3337 -2504 3371 -2488
rect 3595 2488 3629 2504
rect 3595 -2504 3629 -2488
rect 3853 2488 3887 2504
rect 3853 -2504 3887 -2488
rect 4111 2488 4145 2504
rect 4111 -2504 4145 -2488
rect 4369 2488 4403 2504
rect 4369 -2504 4403 -2488
rect -4357 -2581 -4341 -2547
rect -4173 -2581 -4157 -2547
rect -4099 -2581 -4083 -2547
rect -3915 -2581 -3899 -2547
rect -3841 -2581 -3825 -2547
rect -3657 -2581 -3641 -2547
rect -3583 -2581 -3567 -2547
rect -3399 -2581 -3383 -2547
rect -3325 -2581 -3309 -2547
rect -3141 -2581 -3125 -2547
rect -3067 -2581 -3051 -2547
rect -2883 -2581 -2867 -2547
rect -2809 -2581 -2793 -2547
rect -2625 -2581 -2609 -2547
rect -2551 -2581 -2535 -2547
rect -2367 -2581 -2351 -2547
rect -2293 -2581 -2277 -2547
rect -2109 -2581 -2093 -2547
rect -2035 -2581 -2019 -2547
rect -1851 -2581 -1835 -2547
rect -1777 -2581 -1761 -2547
rect -1593 -2581 -1577 -2547
rect -1519 -2581 -1503 -2547
rect -1335 -2581 -1319 -2547
rect -1261 -2581 -1245 -2547
rect -1077 -2581 -1061 -2547
rect -1003 -2581 -987 -2547
rect -819 -2581 -803 -2547
rect -745 -2581 -729 -2547
rect -561 -2581 -545 -2547
rect -487 -2581 -471 -2547
rect -303 -2581 -287 -2547
rect -229 -2581 -213 -2547
rect -45 -2581 -29 -2547
rect 29 -2581 45 -2547
rect 213 -2581 229 -2547
rect 287 -2581 303 -2547
rect 471 -2581 487 -2547
rect 545 -2581 561 -2547
rect 729 -2581 745 -2547
rect 803 -2581 819 -2547
rect 987 -2581 1003 -2547
rect 1061 -2581 1077 -2547
rect 1245 -2581 1261 -2547
rect 1319 -2581 1335 -2547
rect 1503 -2581 1519 -2547
rect 1577 -2581 1593 -2547
rect 1761 -2581 1777 -2547
rect 1835 -2581 1851 -2547
rect 2019 -2581 2035 -2547
rect 2093 -2581 2109 -2547
rect 2277 -2581 2293 -2547
rect 2351 -2581 2367 -2547
rect 2535 -2581 2551 -2547
rect 2609 -2581 2625 -2547
rect 2793 -2581 2809 -2547
rect 2867 -2581 2883 -2547
rect 3051 -2581 3067 -2547
rect 3125 -2581 3141 -2547
rect 3309 -2581 3325 -2547
rect 3383 -2581 3399 -2547
rect 3567 -2581 3583 -2547
rect 3641 -2581 3657 -2547
rect 3825 -2581 3841 -2547
rect 3899 -2581 3915 -2547
rect 4083 -2581 4099 -2547
rect 4157 -2581 4173 -2547
rect 4341 -2581 4357 -2547
rect -4537 -2685 -4503 -2623
rect 4503 -2685 4537 -2623
rect -4537 -2719 -4441 -2685
rect 4441 -2719 4537 -2685
<< viali >>
rect -4341 2547 -4173 2581
rect -4083 2547 -3915 2581
rect -3825 2547 -3657 2581
rect -3567 2547 -3399 2581
rect -3309 2547 -3141 2581
rect -3051 2547 -2883 2581
rect -2793 2547 -2625 2581
rect -2535 2547 -2367 2581
rect -2277 2547 -2109 2581
rect -2019 2547 -1851 2581
rect -1761 2547 -1593 2581
rect -1503 2547 -1335 2581
rect -1245 2547 -1077 2581
rect -987 2547 -819 2581
rect -729 2547 -561 2581
rect -471 2547 -303 2581
rect -213 2547 -45 2581
rect 45 2547 213 2581
rect 303 2547 471 2581
rect 561 2547 729 2581
rect 819 2547 987 2581
rect 1077 2547 1245 2581
rect 1335 2547 1503 2581
rect 1593 2547 1761 2581
rect 1851 2547 2019 2581
rect 2109 2547 2277 2581
rect 2367 2547 2535 2581
rect 2625 2547 2793 2581
rect 2883 2547 3051 2581
rect 3141 2547 3309 2581
rect 3399 2547 3567 2581
rect 3657 2547 3825 2581
rect 3915 2547 4083 2581
rect 4173 2547 4341 2581
rect -4403 -2488 -4369 2488
rect -4145 -2488 -4111 2488
rect -3887 -2488 -3853 2488
rect -3629 -2488 -3595 2488
rect -3371 -2488 -3337 2488
rect -3113 -2488 -3079 2488
rect -2855 -2488 -2821 2488
rect -2597 -2488 -2563 2488
rect -2339 -2488 -2305 2488
rect -2081 -2488 -2047 2488
rect -1823 -2488 -1789 2488
rect -1565 -2488 -1531 2488
rect -1307 -2488 -1273 2488
rect -1049 -2488 -1015 2488
rect -791 -2488 -757 2488
rect -533 -2488 -499 2488
rect -275 -2488 -241 2488
rect -17 -2488 17 2488
rect 241 -2488 275 2488
rect 499 -2488 533 2488
rect 757 -2488 791 2488
rect 1015 -2488 1049 2488
rect 1273 -2488 1307 2488
rect 1531 -2488 1565 2488
rect 1789 -2488 1823 2488
rect 2047 -2488 2081 2488
rect 2305 -2488 2339 2488
rect 2563 -2488 2597 2488
rect 2821 -2488 2855 2488
rect 3079 -2488 3113 2488
rect 3337 -2488 3371 2488
rect 3595 -2488 3629 2488
rect 3853 -2488 3887 2488
rect 4111 -2488 4145 2488
rect 4369 -2488 4403 2488
rect -4341 -2581 -4173 -2547
rect -4083 -2581 -3915 -2547
rect -3825 -2581 -3657 -2547
rect -3567 -2581 -3399 -2547
rect -3309 -2581 -3141 -2547
rect -3051 -2581 -2883 -2547
rect -2793 -2581 -2625 -2547
rect -2535 -2581 -2367 -2547
rect -2277 -2581 -2109 -2547
rect -2019 -2581 -1851 -2547
rect -1761 -2581 -1593 -2547
rect -1503 -2581 -1335 -2547
rect -1245 -2581 -1077 -2547
rect -987 -2581 -819 -2547
rect -729 -2581 -561 -2547
rect -471 -2581 -303 -2547
rect -213 -2581 -45 -2547
rect 45 -2581 213 -2547
rect 303 -2581 471 -2547
rect 561 -2581 729 -2547
rect 819 -2581 987 -2547
rect 1077 -2581 1245 -2547
rect 1335 -2581 1503 -2547
rect 1593 -2581 1761 -2547
rect 1851 -2581 2019 -2547
rect 2109 -2581 2277 -2547
rect 2367 -2581 2535 -2547
rect 2625 -2581 2793 -2547
rect 2883 -2581 3051 -2547
rect 3141 -2581 3309 -2547
rect 3399 -2581 3567 -2547
rect 3657 -2581 3825 -2547
rect 3915 -2581 4083 -2547
rect 4173 -2581 4341 -2547
<< metal1 >>
rect -4353 2581 -4161 2587
rect -4353 2547 -4341 2581
rect -4173 2547 -4161 2581
rect -4353 2541 -4161 2547
rect -4095 2581 -3903 2587
rect -4095 2547 -4083 2581
rect -3915 2547 -3903 2581
rect -4095 2541 -3903 2547
rect -3837 2581 -3645 2587
rect -3837 2547 -3825 2581
rect -3657 2547 -3645 2581
rect -3837 2541 -3645 2547
rect -3579 2581 -3387 2587
rect -3579 2547 -3567 2581
rect -3399 2547 -3387 2581
rect -3579 2541 -3387 2547
rect -3321 2581 -3129 2587
rect -3321 2547 -3309 2581
rect -3141 2547 -3129 2581
rect -3321 2541 -3129 2547
rect -3063 2581 -2871 2587
rect -3063 2547 -3051 2581
rect -2883 2547 -2871 2581
rect -3063 2541 -2871 2547
rect -2805 2581 -2613 2587
rect -2805 2547 -2793 2581
rect -2625 2547 -2613 2581
rect -2805 2541 -2613 2547
rect -2547 2581 -2355 2587
rect -2547 2547 -2535 2581
rect -2367 2547 -2355 2581
rect -2547 2541 -2355 2547
rect -2289 2581 -2097 2587
rect -2289 2547 -2277 2581
rect -2109 2547 -2097 2581
rect -2289 2541 -2097 2547
rect -2031 2581 -1839 2587
rect -2031 2547 -2019 2581
rect -1851 2547 -1839 2581
rect -2031 2541 -1839 2547
rect -1773 2581 -1581 2587
rect -1773 2547 -1761 2581
rect -1593 2547 -1581 2581
rect -1773 2541 -1581 2547
rect -1515 2581 -1323 2587
rect -1515 2547 -1503 2581
rect -1335 2547 -1323 2581
rect -1515 2541 -1323 2547
rect -1257 2581 -1065 2587
rect -1257 2547 -1245 2581
rect -1077 2547 -1065 2581
rect -1257 2541 -1065 2547
rect -999 2581 -807 2587
rect -999 2547 -987 2581
rect -819 2547 -807 2581
rect -999 2541 -807 2547
rect -741 2581 -549 2587
rect -741 2547 -729 2581
rect -561 2547 -549 2581
rect -741 2541 -549 2547
rect -483 2581 -291 2587
rect -483 2547 -471 2581
rect -303 2547 -291 2581
rect -483 2541 -291 2547
rect -225 2581 -33 2587
rect -225 2547 -213 2581
rect -45 2547 -33 2581
rect -225 2541 -33 2547
rect 33 2581 225 2587
rect 33 2547 45 2581
rect 213 2547 225 2581
rect 33 2541 225 2547
rect 291 2581 483 2587
rect 291 2547 303 2581
rect 471 2547 483 2581
rect 291 2541 483 2547
rect 549 2581 741 2587
rect 549 2547 561 2581
rect 729 2547 741 2581
rect 549 2541 741 2547
rect 807 2581 999 2587
rect 807 2547 819 2581
rect 987 2547 999 2581
rect 807 2541 999 2547
rect 1065 2581 1257 2587
rect 1065 2547 1077 2581
rect 1245 2547 1257 2581
rect 1065 2541 1257 2547
rect 1323 2581 1515 2587
rect 1323 2547 1335 2581
rect 1503 2547 1515 2581
rect 1323 2541 1515 2547
rect 1581 2581 1773 2587
rect 1581 2547 1593 2581
rect 1761 2547 1773 2581
rect 1581 2541 1773 2547
rect 1839 2581 2031 2587
rect 1839 2547 1851 2581
rect 2019 2547 2031 2581
rect 1839 2541 2031 2547
rect 2097 2581 2289 2587
rect 2097 2547 2109 2581
rect 2277 2547 2289 2581
rect 2097 2541 2289 2547
rect 2355 2581 2547 2587
rect 2355 2547 2367 2581
rect 2535 2547 2547 2581
rect 2355 2541 2547 2547
rect 2613 2581 2805 2587
rect 2613 2547 2625 2581
rect 2793 2547 2805 2581
rect 2613 2541 2805 2547
rect 2871 2581 3063 2587
rect 2871 2547 2883 2581
rect 3051 2547 3063 2581
rect 2871 2541 3063 2547
rect 3129 2581 3321 2587
rect 3129 2547 3141 2581
rect 3309 2547 3321 2581
rect 3129 2541 3321 2547
rect 3387 2581 3579 2587
rect 3387 2547 3399 2581
rect 3567 2547 3579 2581
rect 3387 2541 3579 2547
rect 3645 2581 3837 2587
rect 3645 2547 3657 2581
rect 3825 2547 3837 2581
rect 3645 2541 3837 2547
rect 3903 2581 4095 2587
rect 3903 2547 3915 2581
rect 4083 2547 4095 2581
rect 3903 2541 4095 2547
rect 4161 2581 4353 2587
rect 4161 2547 4173 2581
rect 4341 2547 4353 2581
rect 4161 2541 4353 2547
rect -4409 2488 -4363 2500
rect -4409 -2488 -4403 2488
rect -4369 -2488 -4363 2488
rect -4409 -2500 -4363 -2488
rect -4151 2488 -4105 2500
rect -4151 -2488 -4145 2488
rect -4111 -2488 -4105 2488
rect -4151 -2500 -4105 -2488
rect -3893 2488 -3847 2500
rect -3893 -2488 -3887 2488
rect -3853 -2488 -3847 2488
rect -3893 -2500 -3847 -2488
rect -3635 2488 -3589 2500
rect -3635 -2488 -3629 2488
rect -3595 -2488 -3589 2488
rect -3635 -2500 -3589 -2488
rect -3377 2488 -3331 2500
rect -3377 -2488 -3371 2488
rect -3337 -2488 -3331 2488
rect -3377 -2500 -3331 -2488
rect -3119 2488 -3073 2500
rect -3119 -2488 -3113 2488
rect -3079 -2488 -3073 2488
rect -3119 -2500 -3073 -2488
rect -2861 2488 -2815 2500
rect -2861 -2488 -2855 2488
rect -2821 -2488 -2815 2488
rect -2861 -2500 -2815 -2488
rect -2603 2488 -2557 2500
rect -2603 -2488 -2597 2488
rect -2563 -2488 -2557 2488
rect -2603 -2500 -2557 -2488
rect -2345 2488 -2299 2500
rect -2345 -2488 -2339 2488
rect -2305 -2488 -2299 2488
rect -2345 -2500 -2299 -2488
rect -2087 2488 -2041 2500
rect -2087 -2488 -2081 2488
rect -2047 -2488 -2041 2488
rect -2087 -2500 -2041 -2488
rect -1829 2488 -1783 2500
rect -1829 -2488 -1823 2488
rect -1789 -2488 -1783 2488
rect -1829 -2500 -1783 -2488
rect -1571 2488 -1525 2500
rect -1571 -2488 -1565 2488
rect -1531 -2488 -1525 2488
rect -1571 -2500 -1525 -2488
rect -1313 2488 -1267 2500
rect -1313 -2488 -1307 2488
rect -1273 -2488 -1267 2488
rect -1313 -2500 -1267 -2488
rect -1055 2488 -1009 2500
rect -1055 -2488 -1049 2488
rect -1015 -2488 -1009 2488
rect -1055 -2500 -1009 -2488
rect -797 2488 -751 2500
rect -797 -2488 -791 2488
rect -757 -2488 -751 2488
rect -797 -2500 -751 -2488
rect -539 2488 -493 2500
rect -539 -2488 -533 2488
rect -499 -2488 -493 2488
rect -539 -2500 -493 -2488
rect -281 2488 -235 2500
rect -281 -2488 -275 2488
rect -241 -2488 -235 2488
rect -281 -2500 -235 -2488
rect -23 2488 23 2500
rect -23 -2488 -17 2488
rect 17 -2488 23 2488
rect -23 -2500 23 -2488
rect 235 2488 281 2500
rect 235 -2488 241 2488
rect 275 -2488 281 2488
rect 235 -2500 281 -2488
rect 493 2488 539 2500
rect 493 -2488 499 2488
rect 533 -2488 539 2488
rect 493 -2500 539 -2488
rect 751 2488 797 2500
rect 751 -2488 757 2488
rect 791 -2488 797 2488
rect 751 -2500 797 -2488
rect 1009 2488 1055 2500
rect 1009 -2488 1015 2488
rect 1049 -2488 1055 2488
rect 1009 -2500 1055 -2488
rect 1267 2488 1313 2500
rect 1267 -2488 1273 2488
rect 1307 -2488 1313 2488
rect 1267 -2500 1313 -2488
rect 1525 2488 1571 2500
rect 1525 -2488 1531 2488
rect 1565 -2488 1571 2488
rect 1525 -2500 1571 -2488
rect 1783 2488 1829 2500
rect 1783 -2488 1789 2488
rect 1823 -2488 1829 2488
rect 1783 -2500 1829 -2488
rect 2041 2488 2087 2500
rect 2041 -2488 2047 2488
rect 2081 -2488 2087 2488
rect 2041 -2500 2087 -2488
rect 2299 2488 2345 2500
rect 2299 -2488 2305 2488
rect 2339 -2488 2345 2488
rect 2299 -2500 2345 -2488
rect 2557 2488 2603 2500
rect 2557 -2488 2563 2488
rect 2597 -2488 2603 2488
rect 2557 -2500 2603 -2488
rect 2815 2488 2861 2500
rect 2815 -2488 2821 2488
rect 2855 -2488 2861 2488
rect 2815 -2500 2861 -2488
rect 3073 2488 3119 2500
rect 3073 -2488 3079 2488
rect 3113 -2488 3119 2488
rect 3073 -2500 3119 -2488
rect 3331 2488 3377 2500
rect 3331 -2488 3337 2488
rect 3371 -2488 3377 2488
rect 3331 -2500 3377 -2488
rect 3589 2488 3635 2500
rect 3589 -2488 3595 2488
rect 3629 -2488 3635 2488
rect 3589 -2500 3635 -2488
rect 3847 2488 3893 2500
rect 3847 -2488 3853 2488
rect 3887 -2488 3893 2488
rect 3847 -2500 3893 -2488
rect 4105 2488 4151 2500
rect 4105 -2488 4111 2488
rect 4145 -2488 4151 2488
rect 4105 -2500 4151 -2488
rect 4363 2488 4409 2500
rect 4363 -2488 4369 2488
rect 4403 -2488 4409 2488
rect 4363 -2500 4409 -2488
rect -4353 -2547 -4161 -2541
rect -4353 -2581 -4341 -2547
rect -4173 -2581 -4161 -2547
rect -4353 -2587 -4161 -2581
rect -4095 -2547 -3903 -2541
rect -4095 -2581 -4083 -2547
rect -3915 -2581 -3903 -2547
rect -4095 -2587 -3903 -2581
rect -3837 -2547 -3645 -2541
rect -3837 -2581 -3825 -2547
rect -3657 -2581 -3645 -2547
rect -3837 -2587 -3645 -2581
rect -3579 -2547 -3387 -2541
rect -3579 -2581 -3567 -2547
rect -3399 -2581 -3387 -2547
rect -3579 -2587 -3387 -2581
rect -3321 -2547 -3129 -2541
rect -3321 -2581 -3309 -2547
rect -3141 -2581 -3129 -2547
rect -3321 -2587 -3129 -2581
rect -3063 -2547 -2871 -2541
rect -3063 -2581 -3051 -2547
rect -2883 -2581 -2871 -2547
rect -3063 -2587 -2871 -2581
rect -2805 -2547 -2613 -2541
rect -2805 -2581 -2793 -2547
rect -2625 -2581 -2613 -2547
rect -2805 -2587 -2613 -2581
rect -2547 -2547 -2355 -2541
rect -2547 -2581 -2535 -2547
rect -2367 -2581 -2355 -2547
rect -2547 -2587 -2355 -2581
rect -2289 -2547 -2097 -2541
rect -2289 -2581 -2277 -2547
rect -2109 -2581 -2097 -2547
rect -2289 -2587 -2097 -2581
rect -2031 -2547 -1839 -2541
rect -2031 -2581 -2019 -2547
rect -1851 -2581 -1839 -2547
rect -2031 -2587 -1839 -2581
rect -1773 -2547 -1581 -2541
rect -1773 -2581 -1761 -2547
rect -1593 -2581 -1581 -2547
rect -1773 -2587 -1581 -2581
rect -1515 -2547 -1323 -2541
rect -1515 -2581 -1503 -2547
rect -1335 -2581 -1323 -2547
rect -1515 -2587 -1323 -2581
rect -1257 -2547 -1065 -2541
rect -1257 -2581 -1245 -2547
rect -1077 -2581 -1065 -2547
rect -1257 -2587 -1065 -2581
rect -999 -2547 -807 -2541
rect -999 -2581 -987 -2547
rect -819 -2581 -807 -2547
rect -999 -2587 -807 -2581
rect -741 -2547 -549 -2541
rect -741 -2581 -729 -2547
rect -561 -2581 -549 -2547
rect -741 -2587 -549 -2581
rect -483 -2547 -291 -2541
rect -483 -2581 -471 -2547
rect -303 -2581 -291 -2547
rect -483 -2587 -291 -2581
rect -225 -2547 -33 -2541
rect -225 -2581 -213 -2547
rect -45 -2581 -33 -2547
rect -225 -2587 -33 -2581
rect 33 -2547 225 -2541
rect 33 -2581 45 -2547
rect 213 -2581 225 -2547
rect 33 -2587 225 -2581
rect 291 -2547 483 -2541
rect 291 -2581 303 -2547
rect 471 -2581 483 -2547
rect 291 -2587 483 -2581
rect 549 -2547 741 -2541
rect 549 -2581 561 -2547
rect 729 -2581 741 -2547
rect 549 -2587 741 -2581
rect 807 -2547 999 -2541
rect 807 -2581 819 -2547
rect 987 -2581 999 -2547
rect 807 -2587 999 -2581
rect 1065 -2547 1257 -2541
rect 1065 -2581 1077 -2547
rect 1245 -2581 1257 -2547
rect 1065 -2587 1257 -2581
rect 1323 -2547 1515 -2541
rect 1323 -2581 1335 -2547
rect 1503 -2581 1515 -2547
rect 1323 -2587 1515 -2581
rect 1581 -2547 1773 -2541
rect 1581 -2581 1593 -2547
rect 1761 -2581 1773 -2547
rect 1581 -2587 1773 -2581
rect 1839 -2547 2031 -2541
rect 1839 -2581 1851 -2547
rect 2019 -2581 2031 -2547
rect 1839 -2587 2031 -2581
rect 2097 -2547 2289 -2541
rect 2097 -2581 2109 -2547
rect 2277 -2581 2289 -2547
rect 2097 -2587 2289 -2581
rect 2355 -2547 2547 -2541
rect 2355 -2581 2367 -2547
rect 2535 -2581 2547 -2547
rect 2355 -2587 2547 -2581
rect 2613 -2547 2805 -2541
rect 2613 -2581 2625 -2547
rect 2793 -2581 2805 -2547
rect 2613 -2587 2805 -2581
rect 2871 -2547 3063 -2541
rect 2871 -2581 2883 -2547
rect 3051 -2581 3063 -2547
rect 2871 -2587 3063 -2581
rect 3129 -2547 3321 -2541
rect 3129 -2581 3141 -2547
rect 3309 -2581 3321 -2547
rect 3129 -2587 3321 -2581
rect 3387 -2547 3579 -2541
rect 3387 -2581 3399 -2547
rect 3567 -2581 3579 -2547
rect 3387 -2587 3579 -2581
rect 3645 -2547 3837 -2541
rect 3645 -2581 3657 -2547
rect 3825 -2581 3837 -2547
rect 3645 -2587 3837 -2581
rect 3903 -2547 4095 -2541
rect 3903 -2581 3915 -2547
rect 4083 -2581 4095 -2547
rect 3903 -2587 4095 -2581
rect 4161 -2547 4353 -2541
rect 4161 -2581 4173 -2547
rect 4341 -2581 4353 -2547
rect 4161 -2587 4353 -2581
<< properties >>
string FIXED_BBOX -4520 -2702 4520 2702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 25 l 1 m 1 nf 34 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713393126
<< nwell >>
rect -1906 -717 1906 717
<< mvpmos >>
rect -1648 -420 -1448 420
rect -1390 -420 -1190 420
rect -1132 -420 -932 420
rect -874 -420 -674 420
rect -616 -420 -416 420
rect -358 -420 -158 420
rect -100 -420 100 420
rect 158 -420 358 420
rect 416 -420 616 420
rect 674 -420 874 420
rect 932 -420 1132 420
rect 1190 -420 1390 420
rect 1448 -420 1648 420
<< mvpdiff >>
rect -1706 408 -1648 420
rect -1706 -408 -1694 408
rect -1660 -408 -1648 408
rect -1706 -420 -1648 -408
rect -1448 408 -1390 420
rect -1448 -408 -1436 408
rect -1402 -408 -1390 408
rect -1448 -420 -1390 -408
rect -1190 408 -1132 420
rect -1190 -408 -1178 408
rect -1144 -408 -1132 408
rect -1190 -420 -1132 -408
rect -932 408 -874 420
rect -932 -408 -920 408
rect -886 -408 -874 408
rect -932 -420 -874 -408
rect -674 408 -616 420
rect -674 -408 -662 408
rect -628 -408 -616 408
rect -674 -420 -616 -408
rect -416 408 -358 420
rect -416 -408 -404 408
rect -370 -408 -358 408
rect -416 -420 -358 -408
rect -158 408 -100 420
rect -158 -408 -146 408
rect -112 -408 -100 408
rect -158 -420 -100 -408
rect 100 408 158 420
rect 100 -408 112 408
rect 146 -408 158 408
rect 100 -420 158 -408
rect 358 408 416 420
rect 358 -408 370 408
rect 404 -408 416 408
rect 358 -420 416 -408
rect 616 408 674 420
rect 616 -408 628 408
rect 662 -408 674 408
rect 616 -420 674 -408
rect 874 408 932 420
rect 874 -408 886 408
rect 920 -408 932 408
rect 874 -420 932 -408
rect 1132 408 1190 420
rect 1132 -408 1144 408
rect 1178 -408 1190 408
rect 1132 -420 1190 -408
rect 1390 408 1448 420
rect 1390 -408 1402 408
rect 1436 -408 1448 408
rect 1390 -420 1448 -408
rect 1648 408 1706 420
rect 1648 -408 1660 408
rect 1694 -408 1706 408
rect 1648 -420 1706 -408
<< mvpdiffc >>
rect -1694 -408 -1660 408
rect -1436 -408 -1402 408
rect -1178 -408 -1144 408
rect -920 -408 -886 408
rect -662 -408 -628 408
rect -404 -408 -370 408
rect -146 -408 -112 408
rect 112 -408 146 408
rect 370 -408 404 408
rect 628 -408 662 408
rect 886 -408 920 408
rect 1144 -408 1178 408
rect 1402 -408 1436 408
rect 1660 -408 1694 408
<< mvnsubdiff >>
rect -1840 639 1840 651
rect -1840 605 -1732 639
rect 1732 605 1840 639
rect -1840 593 1840 605
rect -1840 543 -1782 593
rect -1840 -543 -1828 543
rect -1794 -543 -1782 543
rect 1782 543 1840 593
rect -1840 -593 -1782 -543
rect 1782 -543 1794 543
rect 1828 -543 1840 543
rect 1782 -593 1840 -543
rect -1840 -605 1840 -593
rect -1840 -639 -1732 -605
rect 1732 -639 1840 -605
rect -1840 -651 1840 -639
<< mvnsubdiffcont >>
rect -1732 605 1732 639
rect -1828 -543 -1794 543
rect 1794 -543 1828 543
rect -1732 -639 1732 -605
<< poly >>
rect -1614 501 -1482 517
rect -1614 484 -1598 501
rect -1648 467 -1598 484
rect -1498 484 -1482 501
rect -1356 501 -1224 517
rect -1356 484 -1340 501
rect -1498 467 -1448 484
rect -1648 420 -1448 467
rect -1390 467 -1340 484
rect -1240 484 -1224 501
rect -1098 501 -966 517
rect -1098 484 -1082 501
rect -1240 467 -1190 484
rect -1390 420 -1190 467
rect -1132 467 -1082 484
rect -982 484 -966 501
rect -840 501 -708 517
rect -840 484 -824 501
rect -982 467 -932 484
rect -1132 420 -932 467
rect -874 467 -824 484
rect -724 484 -708 501
rect -582 501 -450 517
rect -582 484 -566 501
rect -724 467 -674 484
rect -874 420 -674 467
rect -616 467 -566 484
rect -466 484 -450 501
rect -324 501 -192 517
rect -324 484 -308 501
rect -466 467 -416 484
rect -616 420 -416 467
rect -358 467 -308 484
rect -208 484 -192 501
rect -66 501 66 517
rect -66 484 -50 501
rect -208 467 -158 484
rect -358 420 -158 467
rect -100 467 -50 484
rect 50 484 66 501
rect 192 501 324 517
rect 192 484 208 501
rect 50 467 100 484
rect -100 420 100 467
rect 158 467 208 484
rect 308 484 324 501
rect 450 501 582 517
rect 450 484 466 501
rect 308 467 358 484
rect 158 420 358 467
rect 416 467 466 484
rect 566 484 582 501
rect 708 501 840 517
rect 708 484 724 501
rect 566 467 616 484
rect 416 420 616 467
rect 674 467 724 484
rect 824 484 840 501
rect 966 501 1098 517
rect 966 484 982 501
rect 824 467 874 484
rect 674 420 874 467
rect 932 467 982 484
rect 1082 484 1098 501
rect 1224 501 1356 517
rect 1224 484 1240 501
rect 1082 467 1132 484
rect 932 420 1132 467
rect 1190 467 1240 484
rect 1340 484 1356 501
rect 1482 501 1614 517
rect 1482 484 1498 501
rect 1340 467 1390 484
rect 1190 420 1390 467
rect 1448 467 1498 484
rect 1598 484 1614 501
rect 1598 467 1648 484
rect 1448 420 1648 467
rect -1648 -467 -1448 -420
rect -1648 -484 -1598 -467
rect -1614 -501 -1598 -484
rect -1498 -484 -1448 -467
rect -1390 -467 -1190 -420
rect -1390 -484 -1340 -467
rect -1498 -501 -1482 -484
rect -1614 -517 -1482 -501
rect -1356 -501 -1340 -484
rect -1240 -484 -1190 -467
rect -1132 -467 -932 -420
rect -1132 -484 -1082 -467
rect -1240 -501 -1224 -484
rect -1356 -517 -1224 -501
rect -1098 -501 -1082 -484
rect -982 -484 -932 -467
rect -874 -467 -674 -420
rect -874 -484 -824 -467
rect -982 -501 -966 -484
rect -1098 -517 -966 -501
rect -840 -501 -824 -484
rect -724 -484 -674 -467
rect -616 -467 -416 -420
rect -616 -484 -566 -467
rect -724 -501 -708 -484
rect -840 -517 -708 -501
rect -582 -501 -566 -484
rect -466 -484 -416 -467
rect -358 -467 -158 -420
rect -358 -484 -308 -467
rect -466 -501 -450 -484
rect -582 -517 -450 -501
rect -324 -501 -308 -484
rect -208 -484 -158 -467
rect -100 -467 100 -420
rect -100 -484 -50 -467
rect -208 -501 -192 -484
rect -324 -517 -192 -501
rect -66 -501 -50 -484
rect 50 -484 100 -467
rect 158 -467 358 -420
rect 158 -484 208 -467
rect 50 -501 66 -484
rect -66 -517 66 -501
rect 192 -501 208 -484
rect 308 -484 358 -467
rect 416 -467 616 -420
rect 416 -484 466 -467
rect 308 -501 324 -484
rect 192 -517 324 -501
rect 450 -501 466 -484
rect 566 -484 616 -467
rect 674 -467 874 -420
rect 674 -484 724 -467
rect 566 -501 582 -484
rect 450 -517 582 -501
rect 708 -501 724 -484
rect 824 -484 874 -467
rect 932 -467 1132 -420
rect 932 -484 982 -467
rect 824 -501 840 -484
rect 708 -517 840 -501
rect 966 -501 982 -484
rect 1082 -484 1132 -467
rect 1190 -467 1390 -420
rect 1190 -484 1240 -467
rect 1082 -501 1098 -484
rect 966 -517 1098 -501
rect 1224 -501 1240 -484
rect 1340 -484 1390 -467
rect 1448 -467 1648 -420
rect 1448 -484 1498 -467
rect 1340 -501 1356 -484
rect 1224 -517 1356 -501
rect 1482 -501 1498 -484
rect 1598 -484 1648 -467
rect 1598 -501 1614 -484
rect 1482 -517 1614 -501
<< polycont >>
rect -1598 467 -1498 501
rect -1340 467 -1240 501
rect -1082 467 -982 501
rect -824 467 -724 501
rect -566 467 -466 501
rect -308 467 -208 501
rect -50 467 50 501
rect 208 467 308 501
rect 466 467 566 501
rect 724 467 824 501
rect 982 467 1082 501
rect 1240 467 1340 501
rect 1498 467 1598 501
rect -1598 -501 -1498 -467
rect -1340 -501 -1240 -467
rect -1082 -501 -982 -467
rect -824 -501 -724 -467
rect -566 -501 -466 -467
rect -308 -501 -208 -467
rect -50 -501 50 -467
rect 208 -501 308 -467
rect 466 -501 566 -467
rect 724 -501 824 -467
rect 982 -501 1082 -467
rect 1240 -501 1340 -467
rect 1498 -501 1598 -467
<< locali >>
rect -1828 605 -1732 639
rect 1732 605 1828 639
rect -1828 543 -1794 605
rect 1794 543 1828 605
rect -1614 467 -1598 501
rect -1498 467 -1482 501
rect -1356 467 -1340 501
rect -1240 467 -1224 501
rect -1098 467 -1082 501
rect -982 467 -966 501
rect -840 467 -824 501
rect -724 467 -708 501
rect -582 467 -566 501
rect -466 467 -450 501
rect -324 467 -308 501
rect -208 467 -192 501
rect -66 467 -50 501
rect 50 467 66 501
rect 192 467 208 501
rect 308 467 324 501
rect 450 467 466 501
rect 566 467 582 501
rect 708 467 724 501
rect 824 467 840 501
rect 966 467 982 501
rect 1082 467 1098 501
rect 1224 467 1240 501
rect 1340 467 1356 501
rect 1482 467 1498 501
rect 1598 467 1614 501
rect -1694 408 -1660 424
rect -1694 -424 -1660 -408
rect -1436 408 -1402 424
rect -1436 -424 -1402 -408
rect -1178 408 -1144 424
rect -1178 -424 -1144 -408
rect -920 408 -886 424
rect -920 -424 -886 -408
rect -662 408 -628 424
rect -662 -424 -628 -408
rect -404 408 -370 424
rect -404 -424 -370 -408
rect -146 408 -112 424
rect -146 -424 -112 -408
rect 112 408 146 424
rect 112 -424 146 -408
rect 370 408 404 424
rect 370 -424 404 -408
rect 628 408 662 424
rect 628 -424 662 -408
rect 886 408 920 424
rect 886 -424 920 -408
rect 1144 408 1178 424
rect 1144 -424 1178 -408
rect 1402 408 1436 424
rect 1402 -424 1436 -408
rect 1660 408 1694 424
rect 1660 -424 1694 -408
rect -1614 -501 -1598 -467
rect -1498 -501 -1482 -467
rect -1356 -501 -1340 -467
rect -1240 -501 -1224 -467
rect -1098 -501 -1082 -467
rect -982 -501 -966 -467
rect -840 -501 -824 -467
rect -724 -501 -708 -467
rect -582 -501 -566 -467
rect -466 -501 -450 -467
rect -324 -501 -308 -467
rect -208 -501 -192 -467
rect -66 -501 -50 -467
rect 50 -501 66 -467
rect 192 -501 208 -467
rect 308 -501 324 -467
rect 450 -501 466 -467
rect 566 -501 582 -467
rect 708 -501 724 -467
rect 824 -501 840 -467
rect 966 -501 982 -467
rect 1082 -501 1098 -467
rect 1224 -501 1240 -467
rect 1340 -501 1356 -467
rect 1482 -501 1498 -467
rect 1598 -501 1614 -467
rect -1828 -605 -1794 -543
rect 1794 -605 1828 -543
rect -1828 -639 -1732 -605
rect 1732 -639 1828 -605
<< viali >>
rect -1598 467 -1498 501
rect -1340 467 -1240 501
rect -1082 467 -982 501
rect -824 467 -724 501
rect -566 467 -466 501
rect -308 467 -208 501
rect -50 467 50 501
rect 208 467 308 501
rect 466 467 566 501
rect 724 467 824 501
rect 982 467 1082 501
rect 1240 467 1340 501
rect 1498 467 1598 501
rect -1694 -408 -1660 408
rect -1436 -408 -1402 408
rect -1178 -408 -1144 408
rect -920 -408 -886 408
rect -662 -408 -628 408
rect -404 -408 -370 408
rect -146 -408 -112 408
rect 112 -408 146 408
rect 370 -408 404 408
rect 628 -408 662 408
rect 886 -408 920 408
rect 1144 -408 1178 408
rect 1402 -408 1436 408
rect 1660 -408 1694 408
rect -1598 -501 -1498 -467
rect -1340 -501 -1240 -467
rect -1082 -501 -982 -467
rect -824 -501 -724 -467
rect -566 -501 -466 -467
rect -308 -501 -208 -467
rect -50 -501 50 -467
rect 208 -501 308 -467
rect 466 -501 566 -467
rect 724 -501 824 -467
rect 982 -501 1082 -467
rect 1240 -501 1340 -467
rect 1498 -501 1598 -467
<< metal1 >>
rect -1610 501 -1486 507
rect -1610 467 -1598 501
rect -1498 467 -1486 501
rect -1610 461 -1486 467
rect -1352 501 -1228 507
rect -1352 467 -1340 501
rect -1240 467 -1228 501
rect -1352 461 -1228 467
rect -1094 501 -970 507
rect -1094 467 -1082 501
rect -982 467 -970 501
rect -1094 461 -970 467
rect -836 501 -712 507
rect -836 467 -824 501
rect -724 467 -712 501
rect -836 461 -712 467
rect -578 501 -454 507
rect -578 467 -566 501
rect -466 467 -454 501
rect -578 461 -454 467
rect -320 501 -196 507
rect -320 467 -308 501
rect -208 467 -196 501
rect -320 461 -196 467
rect -62 501 62 507
rect -62 467 -50 501
rect 50 467 62 501
rect -62 461 62 467
rect 196 501 320 507
rect 196 467 208 501
rect 308 467 320 501
rect 196 461 320 467
rect 454 501 578 507
rect 454 467 466 501
rect 566 467 578 501
rect 454 461 578 467
rect 712 501 836 507
rect 712 467 724 501
rect 824 467 836 501
rect 712 461 836 467
rect 970 501 1094 507
rect 970 467 982 501
rect 1082 467 1094 501
rect 970 461 1094 467
rect 1228 501 1352 507
rect 1228 467 1240 501
rect 1340 467 1352 501
rect 1228 461 1352 467
rect 1486 501 1610 507
rect 1486 467 1498 501
rect 1598 467 1610 501
rect 1486 461 1610 467
rect -1700 408 -1654 420
rect -1700 -408 -1694 408
rect -1660 -408 -1654 408
rect -1700 -420 -1654 -408
rect -1442 408 -1396 420
rect -1442 -408 -1436 408
rect -1402 -408 -1396 408
rect -1442 -420 -1396 -408
rect -1184 408 -1138 420
rect -1184 -408 -1178 408
rect -1144 -408 -1138 408
rect -1184 -420 -1138 -408
rect -926 408 -880 420
rect -926 -408 -920 408
rect -886 -408 -880 408
rect -926 -420 -880 -408
rect -668 408 -622 420
rect -668 -408 -662 408
rect -628 -408 -622 408
rect -668 -420 -622 -408
rect -410 408 -364 420
rect -410 -408 -404 408
rect -370 -408 -364 408
rect -410 -420 -364 -408
rect -152 408 -106 420
rect -152 -408 -146 408
rect -112 -408 -106 408
rect -152 -420 -106 -408
rect 106 408 152 420
rect 106 -408 112 408
rect 146 -408 152 408
rect 106 -420 152 -408
rect 364 408 410 420
rect 364 -408 370 408
rect 404 -408 410 408
rect 364 -420 410 -408
rect 622 408 668 420
rect 622 -408 628 408
rect 662 -408 668 408
rect 622 -420 668 -408
rect 880 408 926 420
rect 880 -408 886 408
rect 920 -408 926 408
rect 880 -420 926 -408
rect 1138 408 1184 420
rect 1138 -408 1144 408
rect 1178 -408 1184 408
rect 1138 -420 1184 -408
rect 1396 408 1442 420
rect 1396 -408 1402 408
rect 1436 -408 1442 408
rect 1396 -420 1442 -408
rect 1654 408 1700 420
rect 1654 -408 1660 408
rect 1694 -408 1700 408
rect 1654 -420 1700 -408
rect -1610 -467 -1486 -461
rect -1610 -501 -1598 -467
rect -1498 -501 -1486 -467
rect -1610 -507 -1486 -501
rect -1352 -467 -1228 -461
rect -1352 -501 -1340 -467
rect -1240 -501 -1228 -467
rect -1352 -507 -1228 -501
rect -1094 -467 -970 -461
rect -1094 -501 -1082 -467
rect -982 -501 -970 -467
rect -1094 -507 -970 -501
rect -836 -467 -712 -461
rect -836 -501 -824 -467
rect -724 -501 -712 -467
rect -836 -507 -712 -501
rect -578 -467 -454 -461
rect -578 -501 -566 -467
rect -466 -501 -454 -467
rect -578 -507 -454 -501
rect -320 -467 -196 -461
rect -320 -501 -308 -467
rect -208 -501 -196 -467
rect -320 -507 -196 -501
rect -62 -467 62 -461
rect -62 -501 -50 -467
rect 50 -501 62 -467
rect -62 -507 62 -501
rect 196 -467 320 -461
rect 196 -501 208 -467
rect 308 -501 320 -467
rect 196 -507 320 -501
rect 454 -467 578 -461
rect 454 -501 466 -467
rect 566 -501 578 -467
rect 454 -507 578 -501
rect 712 -467 836 -461
rect 712 -501 724 -467
rect 824 -501 836 -467
rect 712 -507 836 -501
rect 970 -467 1094 -461
rect 970 -501 982 -467
rect 1082 -501 1094 -467
rect 970 -507 1094 -501
rect 1228 -467 1352 -461
rect 1228 -501 1240 -467
rect 1340 -501 1352 -467
rect 1228 -507 1352 -501
rect 1486 -467 1610 -461
rect 1486 -501 1498 -467
rect 1598 -501 1610 -467
rect 1486 -507 1610 -501
<< properties >>
string FIXED_BBOX -1811 -622 1811 622
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.2 l 1 m 1 nf 13 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713660561
<< nwell >>
rect -550 -506 550 506
<< pdiff >>
rect -392 336 -308 348
rect -392 302 -380 336
rect -320 302 -308 336
rect -392 245 -308 302
rect -392 -302 -308 -245
rect -392 -336 -380 -302
rect -320 -336 -308 -302
rect -392 -348 -308 -336
rect -252 336 -168 348
rect -252 302 -240 336
rect -180 302 -168 336
rect -252 245 -168 302
rect -252 -302 -168 -245
rect -252 -336 -240 -302
rect -180 -336 -168 -302
rect -252 -348 -168 -336
rect -112 336 -28 348
rect -112 302 -100 336
rect -40 302 -28 336
rect -112 245 -28 302
rect -112 -302 -28 -245
rect -112 -336 -100 -302
rect -40 -336 -28 -302
rect -112 -348 -28 -336
rect 28 336 112 348
rect 28 302 40 336
rect 100 302 112 336
rect 28 245 112 302
rect 28 -302 112 -245
rect 28 -336 40 -302
rect 100 -336 112 -302
rect 28 -348 112 -336
rect 168 336 252 348
rect 168 302 180 336
rect 240 302 252 336
rect 168 245 252 302
rect 168 -302 252 -245
rect 168 -336 180 -302
rect 240 -336 252 -302
rect 168 -348 252 -336
rect 308 336 392 348
rect 308 302 320 336
rect 380 302 392 336
rect 308 245 392 302
rect 308 -302 392 -245
rect 308 -336 320 -302
rect 380 -336 392 -302
rect 308 -348 392 -336
<< pdiffc >>
rect -380 302 -320 336
rect -380 -336 -320 -302
rect -240 302 -180 336
rect -240 -336 -180 -302
rect -100 302 -40 336
rect -100 -336 -40 -302
rect 40 302 100 336
rect 40 -336 100 -302
rect 180 302 240 336
rect 180 -336 240 -302
rect 320 302 380 336
rect 320 -336 380 -302
<< nsubdiff >>
rect -514 436 -418 470
rect 418 436 514 470
rect -514 374 -480 436
rect 480 374 514 436
rect -514 -436 -480 -374
rect 480 -436 514 -374
rect -514 -470 -418 -436
rect 418 -470 514 -436
<< nsubdiffcont >>
rect -418 436 418 470
rect -514 -374 -480 374
rect 480 -374 514 374
rect -418 -470 418 -436
<< pdiffres >>
rect -392 -245 -308 245
rect -252 -245 -168 245
rect -112 -245 -28 245
rect 28 -245 112 245
rect 168 -245 252 245
rect 308 -245 392 245
<< locali >>
rect -514 436 -418 470
rect 418 436 514 470
rect -514 374 -480 436
rect 480 374 514 436
rect -396 302 -380 336
rect -320 302 -304 336
rect -256 302 -240 336
rect -180 302 -164 336
rect -116 302 -100 336
rect -40 302 -24 336
rect 24 302 40 336
rect 100 302 116 336
rect 164 302 180 336
rect 240 302 256 336
rect 304 302 320 336
rect 380 302 396 336
rect -396 -336 -380 -302
rect -320 -336 -304 -302
rect -256 -336 -240 -302
rect -180 -336 -164 -302
rect -116 -336 -100 -302
rect -40 -336 -24 -302
rect 24 -336 40 -302
rect 100 -336 116 -302
rect 164 -336 180 -302
rect 240 -336 256 -302
rect 304 -336 320 -302
rect 380 -336 396 -302
rect -514 -436 -480 -374
rect 480 -436 514 -374
rect -514 -470 -418 -436
rect 418 -470 514 -436
<< viali >>
rect -380 302 -320 336
rect -240 302 -180 336
rect -100 302 -40 336
rect 40 302 100 336
rect 180 302 240 336
rect 320 302 380 336
rect -380 262 -320 302
rect -240 262 -180 302
rect -100 262 -40 302
rect 40 262 100 302
rect 180 262 240 302
rect 320 262 380 302
rect -380 -302 -320 -262
rect -240 -302 -180 -262
rect -100 -302 -40 -262
rect 40 -302 100 -262
rect 180 -302 240 -262
rect 320 -302 380 -262
rect -380 -336 -320 -302
rect -240 -336 -180 -302
rect -100 -336 -40 -302
rect 40 -336 100 -302
rect 180 -336 240 -302
rect 320 -336 380 -302
<< metal1 >>
rect -386 336 -314 348
rect -386 262 -380 336
rect -320 262 -314 336
rect -386 250 -314 262
rect -246 336 -174 348
rect -246 262 -240 336
rect -180 262 -174 336
rect -246 250 -174 262
rect -106 336 -34 348
rect -106 262 -100 336
rect -40 262 -34 336
rect -106 250 -34 262
rect 34 336 106 348
rect 34 262 40 336
rect 100 262 106 336
rect 34 250 106 262
rect 174 336 246 348
rect 174 262 180 336
rect 240 262 246 336
rect 174 250 246 262
rect 314 336 386 348
rect 314 262 320 336
rect 380 262 386 336
rect 314 250 386 262
rect -386 -262 -314 -250
rect -386 -336 -380 -262
rect -320 -336 -314 -262
rect -386 -348 -314 -336
rect -246 -262 -174 -250
rect -246 -336 -240 -262
rect -180 -336 -174 -262
rect -246 -348 -174 -336
rect -106 -262 -34 -250
rect -106 -336 -100 -262
rect -40 -336 -34 -262
rect -106 -348 -34 -336
rect 34 -262 106 -250
rect 34 -336 40 -262
rect 100 -336 106 -262
rect 34 -348 106 -336
rect 174 -262 246 -250
rect 174 -336 180 -262
rect 240 -336 246 -262
rect 174 -348 246 -336
rect 314 -262 386 -250
rect 314 -336 320 -262
rect 380 -336 386 -262
rect 314 -348 386 -336
<< properties >>
string FIXED_BBOX -497 -453 497 453
string gencell sky130_fd_pr__res_generic_pd
string library sky130
string parameters w 0.42 l 2.45 m 1 nx 6 wmin 0.42 lmin 2.10 rho 197 val 1.206k dummy 0 dw 0.02 term 0.0 sterm 0.0 caplen 0.60 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713233716
<< nwell >>
rect -5131 -1497 5131 1497
<< mvpmos >>
rect -4873 -1200 -4673 1200
rect -4615 -1200 -4415 1200
rect -4357 -1200 -4157 1200
rect -4099 -1200 -3899 1200
rect -3841 -1200 -3641 1200
rect -3583 -1200 -3383 1200
rect -3325 -1200 -3125 1200
rect -3067 -1200 -2867 1200
rect -2809 -1200 -2609 1200
rect -2551 -1200 -2351 1200
rect -2293 -1200 -2093 1200
rect -2035 -1200 -1835 1200
rect -1777 -1200 -1577 1200
rect -1519 -1200 -1319 1200
rect -1261 -1200 -1061 1200
rect -1003 -1200 -803 1200
rect -745 -1200 -545 1200
rect -487 -1200 -287 1200
rect -229 -1200 -29 1200
rect 29 -1200 229 1200
rect 287 -1200 487 1200
rect 545 -1200 745 1200
rect 803 -1200 1003 1200
rect 1061 -1200 1261 1200
rect 1319 -1200 1519 1200
rect 1577 -1200 1777 1200
rect 1835 -1200 2035 1200
rect 2093 -1200 2293 1200
rect 2351 -1200 2551 1200
rect 2609 -1200 2809 1200
rect 2867 -1200 3067 1200
rect 3125 -1200 3325 1200
rect 3383 -1200 3583 1200
rect 3641 -1200 3841 1200
rect 3899 -1200 4099 1200
rect 4157 -1200 4357 1200
rect 4415 -1200 4615 1200
rect 4673 -1200 4873 1200
<< mvpdiff >>
rect -4931 1188 -4873 1200
rect -4931 -1188 -4919 1188
rect -4885 -1188 -4873 1188
rect -4931 -1200 -4873 -1188
rect -4673 1188 -4615 1200
rect -4673 -1188 -4661 1188
rect -4627 -1188 -4615 1188
rect -4673 -1200 -4615 -1188
rect -4415 1188 -4357 1200
rect -4415 -1188 -4403 1188
rect -4369 -1188 -4357 1188
rect -4415 -1200 -4357 -1188
rect -4157 1188 -4099 1200
rect -4157 -1188 -4145 1188
rect -4111 -1188 -4099 1188
rect -4157 -1200 -4099 -1188
rect -3899 1188 -3841 1200
rect -3899 -1188 -3887 1188
rect -3853 -1188 -3841 1188
rect -3899 -1200 -3841 -1188
rect -3641 1188 -3583 1200
rect -3641 -1188 -3629 1188
rect -3595 -1188 -3583 1188
rect -3641 -1200 -3583 -1188
rect -3383 1188 -3325 1200
rect -3383 -1188 -3371 1188
rect -3337 -1188 -3325 1188
rect -3383 -1200 -3325 -1188
rect -3125 1188 -3067 1200
rect -3125 -1188 -3113 1188
rect -3079 -1188 -3067 1188
rect -3125 -1200 -3067 -1188
rect -2867 1188 -2809 1200
rect -2867 -1188 -2855 1188
rect -2821 -1188 -2809 1188
rect -2867 -1200 -2809 -1188
rect -2609 1188 -2551 1200
rect -2609 -1188 -2597 1188
rect -2563 -1188 -2551 1188
rect -2609 -1200 -2551 -1188
rect -2351 1188 -2293 1200
rect -2351 -1188 -2339 1188
rect -2305 -1188 -2293 1188
rect -2351 -1200 -2293 -1188
rect -2093 1188 -2035 1200
rect -2093 -1188 -2081 1188
rect -2047 -1188 -2035 1188
rect -2093 -1200 -2035 -1188
rect -1835 1188 -1777 1200
rect -1835 -1188 -1823 1188
rect -1789 -1188 -1777 1188
rect -1835 -1200 -1777 -1188
rect -1577 1188 -1519 1200
rect -1577 -1188 -1565 1188
rect -1531 -1188 -1519 1188
rect -1577 -1200 -1519 -1188
rect -1319 1188 -1261 1200
rect -1319 -1188 -1307 1188
rect -1273 -1188 -1261 1188
rect -1319 -1200 -1261 -1188
rect -1061 1188 -1003 1200
rect -1061 -1188 -1049 1188
rect -1015 -1188 -1003 1188
rect -1061 -1200 -1003 -1188
rect -803 1188 -745 1200
rect -803 -1188 -791 1188
rect -757 -1188 -745 1188
rect -803 -1200 -745 -1188
rect -545 1188 -487 1200
rect -545 -1188 -533 1188
rect -499 -1188 -487 1188
rect -545 -1200 -487 -1188
rect -287 1188 -229 1200
rect -287 -1188 -275 1188
rect -241 -1188 -229 1188
rect -287 -1200 -229 -1188
rect -29 1188 29 1200
rect -29 -1188 -17 1188
rect 17 -1188 29 1188
rect -29 -1200 29 -1188
rect 229 1188 287 1200
rect 229 -1188 241 1188
rect 275 -1188 287 1188
rect 229 -1200 287 -1188
rect 487 1188 545 1200
rect 487 -1188 499 1188
rect 533 -1188 545 1188
rect 487 -1200 545 -1188
rect 745 1188 803 1200
rect 745 -1188 757 1188
rect 791 -1188 803 1188
rect 745 -1200 803 -1188
rect 1003 1188 1061 1200
rect 1003 -1188 1015 1188
rect 1049 -1188 1061 1188
rect 1003 -1200 1061 -1188
rect 1261 1188 1319 1200
rect 1261 -1188 1273 1188
rect 1307 -1188 1319 1188
rect 1261 -1200 1319 -1188
rect 1519 1188 1577 1200
rect 1519 -1188 1531 1188
rect 1565 -1188 1577 1188
rect 1519 -1200 1577 -1188
rect 1777 1188 1835 1200
rect 1777 -1188 1789 1188
rect 1823 -1188 1835 1188
rect 1777 -1200 1835 -1188
rect 2035 1188 2093 1200
rect 2035 -1188 2047 1188
rect 2081 -1188 2093 1188
rect 2035 -1200 2093 -1188
rect 2293 1188 2351 1200
rect 2293 -1188 2305 1188
rect 2339 -1188 2351 1188
rect 2293 -1200 2351 -1188
rect 2551 1188 2609 1200
rect 2551 -1188 2563 1188
rect 2597 -1188 2609 1188
rect 2551 -1200 2609 -1188
rect 2809 1188 2867 1200
rect 2809 -1188 2821 1188
rect 2855 -1188 2867 1188
rect 2809 -1200 2867 -1188
rect 3067 1188 3125 1200
rect 3067 -1188 3079 1188
rect 3113 -1188 3125 1188
rect 3067 -1200 3125 -1188
rect 3325 1188 3383 1200
rect 3325 -1188 3337 1188
rect 3371 -1188 3383 1188
rect 3325 -1200 3383 -1188
rect 3583 1188 3641 1200
rect 3583 -1188 3595 1188
rect 3629 -1188 3641 1188
rect 3583 -1200 3641 -1188
rect 3841 1188 3899 1200
rect 3841 -1188 3853 1188
rect 3887 -1188 3899 1188
rect 3841 -1200 3899 -1188
rect 4099 1188 4157 1200
rect 4099 -1188 4111 1188
rect 4145 -1188 4157 1188
rect 4099 -1200 4157 -1188
rect 4357 1188 4415 1200
rect 4357 -1188 4369 1188
rect 4403 -1188 4415 1188
rect 4357 -1200 4415 -1188
rect 4615 1188 4673 1200
rect 4615 -1188 4627 1188
rect 4661 -1188 4673 1188
rect 4615 -1200 4673 -1188
rect 4873 1188 4931 1200
rect 4873 -1188 4885 1188
rect 4919 -1188 4931 1188
rect 4873 -1200 4931 -1188
<< mvpdiffc >>
rect -4919 -1188 -4885 1188
rect -4661 -1188 -4627 1188
rect -4403 -1188 -4369 1188
rect -4145 -1188 -4111 1188
rect -3887 -1188 -3853 1188
rect -3629 -1188 -3595 1188
rect -3371 -1188 -3337 1188
rect -3113 -1188 -3079 1188
rect -2855 -1188 -2821 1188
rect -2597 -1188 -2563 1188
rect -2339 -1188 -2305 1188
rect -2081 -1188 -2047 1188
rect -1823 -1188 -1789 1188
rect -1565 -1188 -1531 1188
rect -1307 -1188 -1273 1188
rect -1049 -1188 -1015 1188
rect -791 -1188 -757 1188
rect -533 -1188 -499 1188
rect -275 -1188 -241 1188
rect -17 -1188 17 1188
rect 241 -1188 275 1188
rect 499 -1188 533 1188
rect 757 -1188 791 1188
rect 1015 -1188 1049 1188
rect 1273 -1188 1307 1188
rect 1531 -1188 1565 1188
rect 1789 -1188 1823 1188
rect 2047 -1188 2081 1188
rect 2305 -1188 2339 1188
rect 2563 -1188 2597 1188
rect 2821 -1188 2855 1188
rect 3079 -1188 3113 1188
rect 3337 -1188 3371 1188
rect 3595 -1188 3629 1188
rect 3853 -1188 3887 1188
rect 4111 -1188 4145 1188
rect 4369 -1188 4403 1188
rect 4627 -1188 4661 1188
rect 4885 -1188 4919 1188
<< mvnsubdiff >>
rect -5065 1419 5065 1431
rect -5065 1385 -4957 1419
rect 4957 1385 5065 1419
rect -5065 1373 5065 1385
rect -5065 1323 -5007 1373
rect -5065 -1323 -5053 1323
rect -5019 -1323 -5007 1323
rect 5007 1323 5065 1373
rect -5065 -1373 -5007 -1323
rect 5007 -1323 5019 1323
rect 5053 -1323 5065 1323
rect 5007 -1373 5065 -1323
rect -5065 -1385 5065 -1373
rect -5065 -1419 -4957 -1385
rect 4957 -1419 5065 -1385
rect -5065 -1431 5065 -1419
<< mvnsubdiffcont >>
rect -4957 1385 4957 1419
rect -5053 -1323 -5019 1323
rect 5019 -1323 5053 1323
rect -4957 -1419 4957 -1385
<< poly >>
rect -4873 1281 -4673 1297
rect -4873 1247 -4857 1281
rect -4689 1247 -4673 1281
rect -4873 1200 -4673 1247
rect -4615 1281 -4415 1297
rect -4615 1247 -4599 1281
rect -4431 1247 -4415 1281
rect -4615 1200 -4415 1247
rect -4357 1281 -4157 1297
rect -4357 1247 -4341 1281
rect -4173 1247 -4157 1281
rect -4357 1200 -4157 1247
rect -4099 1281 -3899 1297
rect -4099 1247 -4083 1281
rect -3915 1247 -3899 1281
rect -4099 1200 -3899 1247
rect -3841 1281 -3641 1297
rect -3841 1247 -3825 1281
rect -3657 1247 -3641 1281
rect -3841 1200 -3641 1247
rect -3583 1281 -3383 1297
rect -3583 1247 -3567 1281
rect -3399 1247 -3383 1281
rect -3583 1200 -3383 1247
rect -3325 1281 -3125 1297
rect -3325 1247 -3309 1281
rect -3141 1247 -3125 1281
rect -3325 1200 -3125 1247
rect -3067 1281 -2867 1297
rect -3067 1247 -3051 1281
rect -2883 1247 -2867 1281
rect -3067 1200 -2867 1247
rect -2809 1281 -2609 1297
rect -2809 1247 -2793 1281
rect -2625 1247 -2609 1281
rect -2809 1200 -2609 1247
rect -2551 1281 -2351 1297
rect -2551 1247 -2535 1281
rect -2367 1247 -2351 1281
rect -2551 1200 -2351 1247
rect -2293 1281 -2093 1297
rect -2293 1247 -2277 1281
rect -2109 1247 -2093 1281
rect -2293 1200 -2093 1247
rect -2035 1281 -1835 1297
rect -2035 1247 -2019 1281
rect -1851 1247 -1835 1281
rect -2035 1200 -1835 1247
rect -1777 1281 -1577 1297
rect -1777 1247 -1761 1281
rect -1593 1247 -1577 1281
rect -1777 1200 -1577 1247
rect -1519 1281 -1319 1297
rect -1519 1247 -1503 1281
rect -1335 1247 -1319 1281
rect -1519 1200 -1319 1247
rect -1261 1281 -1061 1297
rect -1261 1247 -1245 1281
rect -1077 1247 -1061 1281
rect -1261 1200 -1061 1247
rect -1003 1281 -803 1297
rect -1003 1247 -987 1281
rect -819 1247 -803 1281
rect -1003 1200 -803 1247
rect -745 1281 -545 1297
rect -745 1247 -729 1281
rect -561 1247 -545 1281
rect -745 1200 -545 1247
rect -487 1281 -287 1297
rect -487 1247 -471 1281
rect -303 1247 -287 1281
rect -487 1200 -287 1247
rect -229 1281 -29 1297
rect -229 1247 -213 1281
rect -45 1247 -29 1281
rect -229 1200 -29 1247
rect 29 1281 229 1297
rect 29 1247 45 1281
rect 213 1247 229 1281
rect 29 1200 229 1247
rect 287 1281 487 1297
rect 287 1247 303 1281
rect 471 1247 487 1281
rect 287 1200 487 1247
rect 545 1281 745 1297
rect 545 1247 561 1281
rect 729 1247 745 1281
rect 545 1200 745 1247
rect 803 1281 1003 1297
rect 803 1247 819 1281
rect 987 1247 1003 1281
rect 803 1200 1003 1247
rect 1061 1281 1261 1297
rect 1061 1247 1077 1281
rect 1245 1247 1261 1281
rect 1061 1200 1261 1247
rect 1319 1281 1519 1297
rect 1319 1247 1335 1281
rect 1503 1247 1519 1281
rect 1319 1200 1519 1247
rect 1577 1281 1777 1297
rect 1577 1247 1593 1281
rect 1761 1247 1777 1281
rect 1577 1200 1777 1247
rect 1835 1281 2035 1297
rect 1835 1247 1851 1281
rect 2019 1247 2035 1281
rect 1835 1200 2035 1247
rect 2093 1281 2293 1297
rect 2093 1247 2109 1281
rect 2277 1247 2293 1281
rect 2093 1200 2293 1247
rect 2351 1281 2551 1297
rect 2351 1247 2367 1281
rect 2535 1247 2551 1281
rect 2351 1200 2551 1247
rect 2609 1281 2809 1297
rect 2609 1247 2625 1281
rect 2793 1247 2809 1281
rect 2609 1200 2809 1247
rect 2867 1281 3067 1297
rect 2867 1247 2883 1281
rect 3051 1247 3067 1281
rect 2867 1200 3067 1247
rect 3125 1281 3325 1297
rect 3125 1247 3141 1281
rect 3309 1247 3325 1281
rect 3125 1200 3325 1247
rect 3383 1281 3583 1297
rect 3383 1247 3399 1281
rect 3567 1247 3583 1281
rect 3383 1200 3583 1247
rect 3641 1281 3841 1297
rect 3641 1247 3657 1281
rect 3825 1247 3841 1281
rect 3641 1200 3841 1247
rect 3899 1281 4099 1297
rect 3899 1247 3915 1281
rect 4083 1247 4099 1281
rect 3899 1200 4099 1247
rect 4157 1281 4357 1297
rect 4157 1247 4173 1281
rect 4341 1247 4357 1281
rect 4157 1200 4357 1247
rect 4415 1281 4615 1297
rect 4415 1247 4431 1281
rect 4599 1247 4615 1281
rect 4415 1200 4615 1247
rect 4673 1281 4873 1297
rect 4673 1247 4689 1281
rect 4857 1247 4873 1281
rect 4673 1200 4873 1247
rect -4873 -1247 -4673 -1200
rect -4873 -1281 -4857 -1247
rect -4689 -1281 -4673 -1247
rect -4873 -1297 -4673 -1281
rect -4615 -1247 -4415 -1200
rect -4615 -1281 -4599 -1247
rect -4431 -1281 -4415 -1247
rect -4615 -1297 -4415 -1281
rect -4357 -1247 -4157 -1200
rect -4357 -1281 -4341 -1247
rect -4173 -1281 -4157 -1247
rect -4357 -1297 -4157 -1281
rect -4099 -1247 -3899 -1200
rect -4099 -1281 -4083 -1247
rect -3915 -1281 -3899 -1247
rect -4099 -1297 -3899 -1281
rect -3841 -1247 -3641 -1200
rect -3841 -1281 -3825 -1247
rect -3657 -1281 -3641 -1247
rect -3841 -1297 -3641 -1281
rect -3583 -1247 -3383 -1200
rect -3583 -1281 -3567 -1247
rect -3399 -1281 -3383 -1247
rect -3583 -1297 -3383 -1281
rect -3325 -1247 -3125 -1200
rect -3325 -1281 -3309 -1247
rect -3141 -1281 -3125 -1247
rect -3325 -1297 -3125 -1281
rect -3067 -1247 -2867 -1200
rect -3067 -1281 -3051 -1247
rect -2883 -1281 -2867 -1247
rect -3067 -1297 -2867 -1281
rect -2809 -1247 -2609 -1200
rect -2809 -1281 -2793 -1247
rect -2625 -1281 -2609 -1247
rect -2809 -1297 -2609 -1281
rect -2551 -1247 -2351 -1200
rect -2551 -1281 -2535 -1247
rect -2367 -1281 -2351 -1247
rect -2551 -1297 -2351 -1281
rect -2293 -1247 -2093 -1200
rect -2293 -1281 -2277 -1247
rect -2109 -1281 -2093 -1247
rect -2293 -1297 -2093 -1281
rect -2035 -1247 -1835 -1200
rect -2035 -1281 -2019 -1247
rect -1851 -1281 -1835 -1247
rect -2035 -1297 -1835 -1281
rect -1777 -1247 -1577 -1200
rect -1777 -1281 -1761 -1247
rect -1593 -1281 -1577 -1247
rect -1777 -1297 -1577 -1281
rect -1519 -1247 -1319 -1200
rect -1519 -1281 -1503 -1247
rect -1335 -1281 -1319 -1247
rect -1519 -1297 -1319 -1281
rect -1261 -1247 -1061 -1200
rect -1261 -1281 -1245 -1247
rect -1077 -1281 -1061 -1247
rect -1261 -1297 -1061 -1281
rect -1003 -1247 -803 -1200
rect -1003 -1281 -987 -1247
rect -819 -1281 -803 -1247
rect -1003 -1297 -803 -1281
rect -745 -1247 -545 -1200
rect -745 -1281 -729 -1247
rect -561 -1281 -545 -1247
rect -745 -1297 -545 -1281
rect -487 -1247 -287 -1200
rect -487 -1281 -471 -1247
rect -303 -1281 -287 -1247
rect -487 -1297 -287 -1281
rect -229 -1247 -29 -1200
rect -229 -1281 -213 -1247
rect -45 -1281 -29 -1247
rect -229 -1297 -29 -1281
rect 29 -1247 229 -1200
rect 29 -1281 45 -1247
rect 213 -1281 229 -1247
rect 29 -1297 229 -1281
rect 287 -1247 487 -1200
rect 287 -1281 303 -1247
rect 471 -1281 487 -1247
rect 287 -1297 487 -1281
rect 545 -1247 745 -1200
rect 545 -1281 561 -1247
rect 729 -1281 745 -1247
rect 545 -1297 745 -1281
rect 803 -1247 1003 -1200
rect 803 -1281 819 -1247
rect 987 -1281 1003 -1247
rect 803 -1297 1003 -1281
rect 1061 -1247 1261 -1200
rect 1061 -1281 1077 -1247
rect 1245 -1281 1261 -1247
rect 1061 -1297 1261 -1281
rect 1319 -1247 1519 -1200
rect 1319 -1281 1335 -1247
rect 1503 -1281 1519 -1247
rect 1319 -1297 1519 -1281
rect 1577 -1247 1777 -1200
rect 1577 -1281 1593 -1247
rect 1761 -1281 1777 -1247
rect 1577 -1297 1777 -1281
rect 1835 -1247 2035 -1200
rect 1835 -1281 1851 -1247
rect 2019 -1281 2035 -1247
rect 1835 -1297 2035 -1281
rect 2093 -1247 2293 -1200
rect 2093 -1281 2109 -1247
rect 2277 -1281 2293 -1247
rect 2093 -1297 2293 -1281
rect 2351 -1247 2551 -1200
rect 2351 -1281 2367 -1247
rect 2535 -1281 2551 -1247
rect 2351 -1297 2551 -1281
rect 2609 -1247 2809 -1200
rect 2609 -1281 2625 -1247
rect 2793 -1281 2809 -1247
rect 2609 -1297 2809 -1281
rect 2867 -1247 3067 -1200
rect 2867 -1281 2883 -1247
rect 3051 -1281 3067 -1247
rect 2867 -1297 3067 -1281
rect 3125 -1247 3325 -1200
rect 3125 -1281 3141 -1247
rect 3309 -1281 3325 -1247
rect 3125 -1297 3325 -1281
rect 3383 -1247 3583 -1200
rect 3383 -1281 3399 -1247
rect 3567 -1281 3583 -1247
rect 3383 -1297 3583 -1281
rect 3641 -1247 3841 -1200
rect 3641 -1281 3657 -1247
rect 3825 -1281 3841 -1247
rect 3641 -1297 3841 -1281
rect 3899 -1247 4099 -1200
rect 3899 -1281 3915 -1247
rect 4083 -1281 4099 -1247
rect 3899 -1297 4099 -1281
rect 4157 -1247 4357 -1200
rect 4157 -1281 4173 -1247
rect 4341 -1281 4357 -1247
rect 4157 -1297 4357 -1281
rect 4415 -1247 4615 -1200
rect 4415 -1281 4431 -1247
rect 4599 -1281 4615 -1247
rect 4415 -1297 4615 -1281
rect 4673 -1247 4873 -1200
rect 4673 -1281 4689 -1247
rect 4857 -1281 4873 -1247
rect 4673 -1297 4873 -1281
<< polycont >>
rect -4857 1247 -4689 1281
rect -4599 1247 -4431 1281
rect -4341 1247 -4173 1281
rect -4083 1247 -3915 1281
rect -3825 1247 -3657 1281
rect -3567 1247 -3399 1281
rect -3309 1247 -3141 1281
rect -3051 1247 -2883 1281
rect -2793 1247 -2625 1281
rect -2535 1247 -2367 1281
rect -2277 1247 -2109 1281
rect -2019 1247 -1851 1281
rect -1761 1247 -1593 1281
rect -1503 1247 -1335 1281
rect -1245 1247 -1077 1281
rect -987 1247 -819 1281
rect -729 1247 -561 1281
rect -471 1247 -303 1281
rect -213 1247 -45 1281
rect 45 1247 213 1281
rect 303 1247 471 1281
rect 561 1247 729 1281
rect 819 1247 987 1281
rect 1077 1247 1245 1281
rect 1335 1247 1503 1281
rect 1593 1247 1761 1281
rect 1851 1247 2019 1281
rect 2109 1247 2277 1281
rect 2367 1247 2535 1281
rect 2625 1247 2793 1281
rect 2883 1247 3051 1281
rect 3141 1247 3309 1281
rect 3399 1247 3567 1281
rect 3657 1247 3825 1281
rect 3915 1247 4083 1281
rect 4173 1247 4341 1281
rect 4431 1247 4599 1281
rect 4689 1247 4857 1281
rect -4857 -1281 -4689 -1247
rect -4599 -1281 -4431 -1247
rect -4341 -1281 -4173 -1247
rect -4083 -1281 -3915 -1247
rect -3825 -1281 -3657 -1247
rect -3567 -1281 -3399 -1247
rect -3309 -1281 -3141 -1247
rect -3051 -1281 -2883 -1247
rect -2793 -1281 -2625 -1247
rect -2535 -1281 -2367 -1247
rect -2277 -1281 -2109 -1247
rect -2019 -1281 -1851 -1247
rect -1761 -1281 -1593 -1247
rect -1503 -1281 -1335 -1247
rect -1245 -1281 -1077 -1247
rect -987 -1281 -819 -1247
rect -729 -1281 -561 -1247
rect -471 -1281 -303 -1247
rect -213 -1281 -45 -1247
rect 45 -1281 213 -1247
rect 303 -1281 471 -1247
rect 561 -1281 729 -1247
rect 819 -1281 987 -1247
rect 1077 -1281 1245 -1247
rect 1335 -1281 1503 -1247
rect 1593 -1281 1761 -1247
rect 1851 -1281 2019 -1247
rect 2109 -1281 2277 -1247
rect 2367 -1281 2535 -1247
rect 2625 -1281 2793 -1247
rect 2883 -1281 3051 -1247
rect 3141 -1281 3309 -1247
rect 3399 -1281 3567 -1247
rect 3657 -1281 3825 -1247
rect 3915 -1281 4083 -1247
rect 4173 -1281 4341 -1247
rect 4431 -1281 4599 -1247
rect 4689 -1281 4857 -1247
<< locali >>
rect -5053 1385 -4957 1419
rect 4957 1385 5053 1419
rect -5053 1323 -5019 1385
rect 5019 1323 5053 1385
rect -4873 1247 -4857 1281
rect -4689 1247 -4673 1281
rect -4615 1247 -4599 1281
rect -4431 1247 -4415 1281
rect -4357 1247 -4341 1281
rect -4173 1247 -4157 1281
rect -4099 1247 -4083 1281
rect -3915 1247 -3899 1281
rect -3841 1247 -3825 1281
rect -3657 1247 -3641 1281
rect -3583 1247 -3567 1281
rect -3399 1247 -3383 1281
rect -3325 1247 -3309 1281
rect -3141 1247 -3125 1281
rect -3067 1247 -3051 1281
rect -2883 1247 -2867 1281
rect -2809 1247 -2793 1281
rect -2625 1247 -2609 1281
rect -2551 1247 -2535 1281
rect -2367 1247 -2351 1281
rect -2293 1247 -2277 1281
rect -2109 1247 -2093 1281
rect -2035 1247 -2019 1281
rect -1851 1247 -1835 1281
rect -1777 1247 -1761 1281
rect -1593 1247 -1577 1281
rect -1519 1247 -1503 1281
rect -1335 1247 -1319 1281
rect -1261 1247 -1245 1281
rect -1077 1247 -1061 1281
rect -1003 1247 -987 1281
rect -819 1247 -803 1281
rect -745 1247 -729 1281
rect -561 1247 -545 1281
rect -487 1247 -471 1281
rect -303 1247 -287 1281
rect -229 1247 -213 1281
rect -45 1247 -29 1281
rect 29 1247 45 1281
rect 213 1247 229 1281
rect 287 1247 303 1281
rect 471 1247 487 1281
rect 545 1247 561 1281
rect 729 1247 745 1281
rect 803 1247 819 1281
rect 987 1247 1003 1281
rect 1061 1247 1077 1281
rect 1245 1247 1261 1281
rect 1319 1247 1335 1281
rect 1503 1247 1519 1281
rect 1577 1247 1593 1281
rect 1761 1247 1777 1281
rect 1835 1247 1851 1281
rect 2019 1247 2035 1281
rect 2093 1247 2109 1281
rect 2277 1247 2293 1281
rect 2351 1247 2367 1281
rect 2535 1247 2551 1281
rect 2609 1247 2625 1281
rect 2793 1247 2809 1281
rect 2867 1247 2883 1281
rect 3051 1247 3067 1281
rect 3125 1247 3141 1281
rect 3309 1247 3325 1281
rect 3383 1247 3399 1281
rect 3567 1247 3583 1281
rect 3641 1247 3657 1281
rect 3825 1247 3841 1281
rect 3899 1247 3915 1281
rect 4083 1247 4099 1281
rect 4157 1247 4173 1281
rect 4341 1247 4357 1281
rect 4415 1247 4431 1281
rect 4599 1247 4615 1281
rect 4673 1247 4689 1281
rect 4857 1247 4873 1281
rect -4919 1188 -4885 1204
rect -4919 -1204 -4885 -1188
rect -4661 1188 -4627 1204
rect -4661 -1204 -4627 -1188
rect -4403 1188 -4369 1204
rect -4403 -1204 -4369 -1188
rect -4145 1188 -4111 1204
rect -4145 -1204 -4111 -1188
rect -3887 1188 -3853 1204
rect -3887 -1204 -3853 -1188
rect -3629 1188 -3595 1204
rect -3629 -1204 -3595 -1188
rect -3371 1188 -3337 1204
rect -3371 -1204 -3337 -1188
rect -3113 1188 -3079 1204
rect -3113 -1204 -3079 -1188
rect -2855 1188 -2821 1204
rect -2855 -1204 -2821 -1188
rect -2597 1188 -2563 1204
rect -2597 -1204 -2563 -1188
rect -2339 1188 -2305 1204
rect -2339 -1204 -2305 -1188
rect -2081 1188 -2047 1204
rect -2081 -1204 -2047 -1188
rect -1823 1188 -1789 1204
rect -1823 -1204 -1789 -1188
rect -1565 1188 -1531 1204
rect -1565 -1204 -1531 -1188
rect -1307 1188 -1273 1204
rect -1307 -1204 -1273 -1188
rect -1049 1188 -1015 1204
rect -1049 -1204 -1015 -1188
rect -791 1188 -757 1204
rect -791 -1204 -757 -1188
rect -533 1188 -499 1204
rect -533 -1204 -499 -1188
rect -275 1188 -241 1204
rect -275 -1204 -241 -1188
rect -17 1188 17 1204
rect -17 -1204 17 -1188
rect 241 1188 275 1204
rect 241 -1204 275 -1188
rect 499 1188 533 1204
rect 499 -1204 533 -1188
rect 757 1188 791 1204
rect 757 -1204 791 -1188
rect 1015 1188 1049 1204
rect 1015 -1204 1049 -1188
rect 1273 1188 1307 1204
rect 1273 -1204 1307 -1188
rect 1531 1188 1565 1204
rect 1531 -1204 1565 -1188
rect 1789 1188 1823 1204
rect 1789 -1204 1823 -1188
rect 2047 1188 2081 1204
rect 2047 -1204 2081 -1188
rect 2305 1188 2339 1204
rect 2305 -1204 2339 -1188
rect 2563 1188 2597 1204
rect 2563 -1204 2597 -1188
rect 2821 1188 2855 1204
rect 2821 -1204 2855 -1188
rect 3079 1188 3113 1204
rect 3079 -1204 3113 -1188
rect 3337 1188 3371 1204
rect 3337 -1204 3371 -1188
rect 3595 1188 3629 1204
rect 3595 -1204 3629 -1188
rect 3853 1188 3887 1204
rect 3853 -1204 3887 -1188
rect 4111 1188 4145 1204
rect 4111 -1204 4145 -1188
rect 4369 1188 4403 1204
rect 4369 -1204 4403 -1188
rect 4627 1188 4661 1204
rect 4627 -1204 4661 -1188
rect 4885 1188 4919 1204
rect 4885 -1204 4919 -1188
rect -4873 -1281 -4857 -1247
rect -4689 -1281 -4673 -1247
rect -4615 -1281 -4599 -1247
rect -4431 -1281 -4415 -1247
rect -4357 -1281 -4341 -1247
rect -4173 -1281 -4157 -1247
rect -4099 -1281 -4083 -1247
rect -3915 -1281 -3899 -1247
rect -3841 -1281 -3825 -1247
rect -3657 -1281 -3641 -1247
rect -3583 -1281 -3567 -1247
rect -3399 -1281 -3383 -1247
rect -3325 -1281 -3309 -1247
rect -3141 -1281 -3125 -1247
rect -3067 -1281 -3051 -1247
rect -2883 -1281 -2867 -1247
rect -2809 -1281 -2793 -1247
rect -2625 -1281 -2609 -1247
rect -2551 -1281 -2535 -1247
rect -2367 -1281 -2351 -1247
rect -2293 -1281 -2277 -1247
rect -2109 -1281 -2093 -1247
rect -2035 -1281 -2019 -1247
rect -1851 -1281 -1835 -1247
rect -1777 -1281 -1761 -1247
rect -1593 -1281 -1577 -1247
rect -1519 -1281 -1503 -1247
rect -1335 -1281 -1319 -1247
rect -1261 -1281 -1245 -1247
rect -1077 -1281 -1061 -1247
rect -1003 -1281 -987 -1247
rect -819 -1281 -803 -1247
rect -745 -1281 -729 -1247
rect -561 -1281 -545 -1247
rect -487 -1281 -471 -1247
rect -303 -1281 -287 -1247
rect -229 -1281 -213 -1247
rect -45 -1281 -29 -1247
rect 29 -1281 45 -1247
rect 213 -1281 229 -1247
rect 287 -1281 303 -1247
rect 471 -1281 487 -1247
rect 545 -1281 561 -1247
rect 729 -1281 745 -1247
rect 803 -1281 819 -1247
rect 987 -1281 1003 -1247
rect 1061 -1281 1077 -1247
rect 1245 -1281 1261 -1247
rect 1319 -1281 1335 -1247
rect 1503 -1281 1519 -1247
rect 1577 -1281 1593 -1247
rect 1761 -1281 1777 -1247
rect 1835 -1281 1851 -1247
rect 2019 -1281 2035 -1247
rect 2093 -1281 2109 -1247
rect 2277 -1281 2293 -1247
rect 2351 -1281 2367 -1247
rect 2535 -1281 2551 -1247
rect 2609 -1281 2625 -1247
rect 2793 -1281 2809 -1247
rect 2867 -1281 2883 -1247
rect 3051 -1281 3067 -1247
rect 3125 -1281 3141 -1247
rect 3309 -1281 3325 -1247
rect 3383 -1281 3399 -1247
rect 3567 -1281 3583 -1247
rect 3641 -1281 3657 -1247
rect 3825 -1281 3841 -1247
rect 3899 -1281 3915 -1247
rect 4083 -1281 4099 -1247
rect 4157 -1281 4173 -1247
rect 4341 -1281 4357 -1247
rect 4415 -1281 4431 -1247
rect 4599 -1281 4615 -1247
rect 4673 -1281 4689 -1247
rect 4857 -1281 4873 -1247
rect -5053 -1385 -5019 -1323
rect 5019 -1385 5053 -1323
rect -5053 -1419 -4957 -1385
rect 4957 -1419 5053 -1385
<< viali >>
rect -4857 1247 -4689 1281
rect -4599 1247 -4431 1281
rect -4341 1247 -4173 1281
rect -4083 1247 -3915 1281
rect -3825 1247 -3657 1281
rect -3567 1247 -3399 1281
rect -3309 1247 -3141 1281
rect -3051 1247 -2883 1281
rect -2793 1247 -2625 1281
rect -2535 1247 -2367 1281
rect -2277 1247 -2109 1281
rect -2019 1247 -1851 1281
rect -1761 1247 -1593 1281
rect -1503 1247 -1335 1281
rect -1245 1247 -1077 1281
rect -987 1247 -819 1281
rect -729 1247 -561 1281
rect -471 1247 -303 1281
rect -213 1247 -45 1281
rect 45 1247 213 1281
rect 303 1247 471 1281
rect 561 1247 729 1281
rect 819 1247 987 1281
rect 1077 1247 1245 1281
rect 1335 1247 1503 1281
rect 1593 1247 1761 1281
rect 1851 1247 2019 1281
rect 2109 1247 2277 1281
rect 2367 1247 2535 1281
rect 2625 1247 2793 1281
rect 2883 1247 3051 1281
rect 3141 1247 3309 1281
rect 3399 1247 3567 1281
rect 3657 1247 3825 1281
rect 3915 1247 4083 1281
rect 4173 1247 4341 1281
rect 4431 1247 4599 1281
rect 4689 1247 4857 1281
rect -4919 -1188 -4885 1188
rect -4661 -1188 -4627 1188
rect -4403 -1188 -4369 1188
rect -4145 -1188 -4111 1188
rect -3887 -1188 -3853 1188
rect -3629 -1188 -3595 1188
rect -3371 -1188 -3337 1188
rect -3113 -1188 -3079 1188
rect -2855 -1188 -2821 1188
rect -2597 -1188 -2563 1188
rect -2339 -1188 -2305 1188
rect -2081 -1188 -2047 1188
rect -1823 -1188 -1789 1188
rect -1565 -1188 -1531 1188
rect -1307 -1188 -1273 1188
rect -1049 -1188 -1015 1188
rect -791 -1188 -757 1188
rect -533 -1188 -499 1188
rect -275 -1188 -241 1188
rect -17 -1188 17 1188
rect 241 -1188 275 1188
rect 499 -1188 533 1188
rect 757 -1188 791 1188
rect 1015 -1188 1049 1188
rect 1273 -1188 1307 1188
rect 1531 -1188 1565 1188
rect 1789 -1188 1823 1188
rect 2047 -1188 2081 1188
rect 2305 -1188 2339 1188
rect 2563 -1188 2597 1188
rect 2821 -1188 2855 1188
rect 3079 -1188 3113 1188
rect 3337 -1188 3371 1188
rect 3595 -1188 3629 1188
rect 3853 -1188 3887 1188
rect 4111 -1188 4145 1188
rect 4369 -1188 4403 1188
rect 4627 -1188 4661 1188
rect 4885 -1188 4919 1188
rect -4857 -1281 -4689 -1247
rect -4599 -1281 -4431 -1247
rect -4341 -1281 -4173 -1247
rect -4083 -1281 -3915 -1247
rect -3825 -1281 -3657 -1247
rect -3567 -1281 -3399 -1247
rect -3309 -1281 -3141 -1247
rect -3051 -1281 -2883 -1247
rect -2793 -1281 -2625 -1247
rect -2535 -1281 -2367 -1247
rect -2277 -1281 -2109 -1247
rect -2019 -1281 -1851 -1247
rect -1761 -1281 -1593 -1247
rect -1503 -1281 -1335 -1247
rect -1245 -1281 -1077 -1247
rect -987 -1281 -819 -1247
rect -729 -1281 -561 -1247
rect -471 -1281 -303 -1247
rect -213 -1281 -45 -1247
rect 45 -1281 213 -1247
rect 303 -1281 471 -1247
rect 561 -1281 729 -1247
rect 819 -1281 987 -1247
rect 1077 -1281 1245 -1247
rect 1335 -1281 1503 -1247
rect 1593 -1281 1761 -1247
rect 1851 -1281 2019 -1247
rect 2109 -1281 2277 -1247
rect 2367 -1281 2535 -1247
rect 2625 -1281 2793 -1247
rect 2883 -1281 3051 -1247
rect 3141 -1281 3309 -1247
rect 3399 -1281 3567 -1247
rect 3657 -1281 3825 -1247
rect 3915 -1281 4083 -1247
rect 4173 -1281 4341 -1247
rect 4431 -1281 4599 -1247
rect 4689 -1281 4857 -1247
<< metal1 >>
rect -4869 1281 -4677 1287
rect -4869 1247 -4857 1281
rect -4689 1247 -4677 1281
rect -4869 1241 -4677 1247
rect -4611 1281 -4419 1287
rect -4611 1247 -4599 1281
rect -4431 1247 -4419 1281
rect -4611 1241 -4419 1247
rect -4353 1281 -4161 1287
rect -4353 1247 -4341 1281
rect -4173 1247 -4161 1281
rect -4353 1241 -4161 1247
rect -4095 1281 -3903 1287
rect -4095 1247 -4083 1281
rect -3915 1247 -3903 1281
rect -4095 1241 -3903 1247
rect -3837 1281 -3645 1287
rect -3837 1247 -3825 1281
rect -3657 1247 -3645 1281
rect -3837 1241 -3645 1247
rect -3579 1281 -3387 1287
rect -3579 1247 -3567 1281
rect -3399 1247 -3387 1281
rect -3579 1241 -3387 1247
rect -3321 1281 -3129 1287
rect -3321 1247 -3309 1281
rect -3141 1247 -3129 1281
rect -3321 1241 -3129 1247
rect -3063 1281 -2871 1287
rect -3063 1247 -3051 1281
rect -2883 1247 -2871 1281
rect -3063 1241 -2871 1247
rect -2805 1281 -2613 1287
rect -2805 1247 -2793 1281
rect -2625 1247 -2613 1281
rect -2805 1241 -2613 1247
rect -2547 1281 -2355 1287
rect -2547 1247 -2535 1281
rect -2367 1247 -2355 1281
rect -2547 1241 -2355 1247
rect -2289 1281 -2097 1287
rect -2289 1247 -2277 1281
rect -2109 1247 -2097 1281
rect -2289 1241 -2097 1247
rect -2031 1281 -1839 1287
rect -2031 1247 -2019 1281
rect -1851 1247 -1839 1281
rect -2031 1241 -1839 1247
rect -1773 1281 -1581 1287
rect -1773 1247 -1761 1281
rect -1593 1247 -1581 1281
rect -1773 1241 -1581 1247
rect -1515 1281 -1323 1287
rect -1515 1247 -1503 1281
rect -1335 1247 -1323 1281
rect -1515 1241 -1323 1247
rect -1257 1281 -1065 1287
rect -1257 1247 -1245 1281
rect -1077 1247 -1065 1281
rect -1257 1241 -1065 1247
rect -999 1281 -807 1287
rect -999 1247 -987 1281
rect -819 1247 -807 1281
rect -999 1241 -807 1247
rect -741 1281 -549 1287
rect -741 1247 -729 1281
rect -561 1247 -549 1281
rect -741 1241 -549 1247
rect -483 1281 -291 1287
rect -483 1247 -471 1281
rect -303 1247 -291 1281
rect -483 1241 -291 1247
rect -225 1281 -33 1287
rect -225 1247 -213 1281
rect -45 1247 -33 1281
rect -225 1241 -33 1247
rect 33 1281 225 1287
rect 33 1247 45 1281
rect 213 1247 225 1281
rect 33 1241 225 1247
rect 291 1281 483 1287
rect 291 1247 303 1281
rect 471 1247 483 1281
rect 291 1241 483 1247
rect 549 1281 741 1287
rect 549 1247 561 1281
rect 729 1247 741 1281
rect 549 1241 741 1247
rect 807 1281 999 1287
rect 807 1247 819 1281
rect 987 1247 999 1281
rect 807 1241 999 1247
rect 1065 1281 1257 1287
rect 1065 1247 1077 1281
rect 1245 1247 1257 1281
rect 1065 1241 1257 1247
rect 1323 1281 1515 1287
rect 1323 1247 1335 1281
rect 1503 1247 1515 1281
rect 1323 1241 1515 1247
rect 1581 1281 1773 1287
rect 1581 1247 1593 1281
rect 1761 1247 1773 1281
rect 1581 1241 1773 1247
rect 1839 1281 2031 1287
rect 1839 1247 1851 1281
rect 2019 1247 2031 1281
rect 1839 1241 2031 1247
rect 2097 1281 2289 1287
rect 2097 1247 2109 1281
rect 2277 1247 2289 1281
rect 2097 1241 2289 1247
rect 2355 1281 2547 1287
rect 2355 1247 2367 1281
rect 2535 1247 2547 1281
rect 2355 1241 2547 1247
rect 2613 1281 2805 1287
rect 2613 1247 2625 1281
rect 2793 1247 2805 1281
rect 2613 1241 2805 1247
rect 2871 1281 3063 1287
rect 2871 1247 2883 1281
rect 3051 1247 3063 1281
rect 2871 1241 3063 1247
rect 3129 1281 3321 1287
rect 3129 1247 3141 1281
rect 3309 1247 3321 1281
rect 3129 1241 3321 1247
rect 3387 1281 3579 1287
rect 3387 1247 3399 1281
rect 3567 1247 3579 1281
rect 3387 1241 3579 1247
rect 3645 1281 3837 1287
rect 3645 1247 3657 1281
rect 3825 1247 3837 1281
rect 3645 1241 3837 1247
rect 3903 1281 4095 1287
rect 3903 1247 3915 1281
rect 4083 1247 4095 1281
rect 3903 1241 4095 1247
rect 4161 1281 4353 1287
rect 4161 1247 4173 1281
rect 4341 1247 4353 1281
rect 4161 1241 4353 1247
rect 4419 1281 4611 1287
rect 4419 1247 4431 1281
rect 4599 1247 4611 1281
rect 4419 1241 4611 1247
rect 4677 1281 4869 1287
rect 4677 1247 4689 1281
rect 4857 1247 4869 1281
rect 4677 1241 4869 1247
rect -4925 1188 -4879 1200
rect -4925 -1188 -4919 1188
rect -4885 -1188 -4879 1188
rect -4925 -1200 -4879 -1188
rect -4667 1188 -4621 1200
rect -4667 -1188 -4661 1188
rect -4627 -1188 -4621 1188
rect -4667 -1200 -4621 -1188
rect -4409 1188 -4363 1200
rect -4409 -1188 -4403 1188
rect -4369 -1188 -4363 1188
rect -4409 -1200 -4363 -1188
rect -4151 1188 -4105 1200
rect -4151 -1188 -4145 1188
rect -4111 -1188 -4105 1188
rect -4151 -1200 -4105 -1188
rect -3893 1188 -3847 1200
rect -3893 -1188 -3887 1188
rect -3853 -1188 -3847 1188
rect -3893 -1200 -3847 -1188
rect -3635 1188 -3589 1200
rect -3635 -1188 -3629 1188
rect -3595 -1188 -3589 1188
rect -3635 -1200 -3589 -1188
rect -3377 1188 -3331 1200
rect -3377 -1188 -3371 1188
rect -3337 -1188 -3331 1188
rect -3377 -1200 -3331 -1188
rect -3119 1188 -3073 1200
rect -3119 -1188 -3113 1188
rect -3079 -1188 -3073 1188
rect -3119 -1200 -3073 -1188
rect -2861 1188 -2815 1200
rect -2861 -1188 -2855 1188
rect -2821 -1188 -2815 1188
rect -2861 -1200 -2815 -1188
rect -2603 1188 -2557 1200
rect -2603 -1188 -2597 1188
rect -2563 -1188 -2557 1188
rect -2603 -1200 -2557 -1188
rect -2345 1188 -2299 1200
rect -2345 -1188 -2339 1188
rect -2305 -1188 -2299 1188
rect -2345 -1200 -2299 -1188
rect -2087 1188 -2041 1200
rect -2087 -1188 -2081 1188
rect -2047 -1188 -2041 1188
rect -2087 -1200 -2041 -1188
rect -1829 1188 -1783 1200
rect -1829 -1188 -1823 1188
rect -1789 -1188 -1783 1188
rect -1829 -1200 -1783 -1188
rect -1571 1188 -1525 1200
rect -1571 -1188 -1565 1188
rect -1531 -1188 -1525 1188
rect -1571 -1200 -1525 -1188
rect -1313 1188 -1267 1200
rect -1313 -1188 -1307 1188
rect -1273 -1188 -1267 1188
rect -1313 -1200 -1267 -1188
rect -1055 1188 -1009 1200
rect -1055 -1188 -1049 1188
rect -1015 -1188 -1009 1188
rect -1055 -1200 -1009 -1188
rect -797 1188 -751 1200
rect -797 -1188 -791 1188
rect -757 -1188 -751 1188
rect -797 -1200 -751 -1188
rect -539 1188 -493 1200
rect -539 -1188 -533 1188
rect -499 -1188 -493 1188
rect -539 -1200 -493 -1188
rect -281 1188 -235 1200
rect -281 -1188 -275 1188
rect -241 -1188 -235 1188
rect -281 -1200 -235 -1188
rect -23 1188 23 1200
rect -23 -1188 -17 1188
rect 17 -1188 23 1188
rect -23 -1200 23 -1188
rect 235 1188 281 1200
rect 235 -1188 241 1188
rect 275 -1188 281 1188
rect 235 -1200 281 -1188
rect 493 1188 539 1200
rect 493 -1188 499 1188
rect 533 -1188 539 1188
rect 493 -1200 539 -1188
rect 751 1188 797 1200
rect 751 -1188 757 1188
rect 791 -1188 797 1188
rect 751 -1200 797 -1188
rect 1009 1188 1055 1200
rect 1009 -1188 1015 1188
rect 1049 -1188 1055 1188
rect 1009 -1200 1055 -1188
rect 1267 1188 1313 1200
rect 1267 -1188 1273 1188
rect 1307 -1188 1313 1188
rect 1267 -1200 1313 -1188
rect 1525 1188 1571 1200
rect 1525 -1188 1531 1188
rect 1565 -1188 1571 1188
rect 1525 -1200 1571 -1188
rect 1783 1188 1829 1200
rect 1783 -1188 1789 1188
rect 1823 -1188 1829 1188
rect 1783 -1200 1829 -1188
rect 2041 1188 2087 1200
rect 2041 -1188 2047 1188
rect 2081 -1188 2087 1188
rect 2041 -1200 2087 -1188
rect 2299 1188 2345 1200
rect 2299 -1188 2305 1188
rect 2339 -1188 2345 1188
rect 2299 -1200 2345 -1188
rect 2557 1188 2603 1200
rect 2557 -1188 2563 1188
rect 2597 -1188 2603 1188
rect 2557 -1200 2603 -1188
rect 2815 1188 2861 1200
rect 2815 -1188 2821 1188
rect 2855 -1188 2861 1188
rect 2815 -1200 2861 -1188
rect 3073 1188 3119 1200
rect 3073 -1188 3079 1188
rect 3113 -1188 3119 1188
rect 3073 -1200 3119 -1188
rect 3331 1188 3377 1200
rect 3331 -1188 3337 1188
rect 3371 -1188 3377 1188
rect 3331 -1200 3377 -1188
rect 3589 1188 3635 1200
rect 3589 -1188 3595 1188
rect 3629 -1188 3635 1188
rect 3589 -1200 3635 -1188
rect 3847 1188 3893 1200
rect 3847 -1188 3853 1188
rect 3887 -1188 3893 1188
rect 3847 -1200 3893 -1188
rect 4105 1188 4151 1200
rect 4105 -1188 4111 1188
rect 4145 -1188 4151 1188
rect 4105 -1200 4151 -1188
rect 4363 1188 4409 1200
rect 4363 -1188 4369 1188
rect 4403 -1188 4409 1188
rect 4363 -1200 4409 -1188
rect 4621 1188 4667 1200
rect 4621 -1188 4627 1188
rect 4661 -1188 4667 1188
rect 4621 -1200 4667 -1188
rect 4879 1188 4925 1200
rect 4879 -1188 4885 1188
rect 4919 -1188 4925 1188
rect 4879 -1200 4925 -1188
rect -4869 -1247 -4677 -1241
rect -4869 -1281 -4857 -1247
rect -4689 -1281 -4677 -1247
rect -4869 -1287 -4677 -1281
rect -4611 -1247 -4419 -1241
rect -4611 -1281 -4599 -1247
rect -4431 -1281 -4419 -1247
rect -4611 -1287 -4419 -1281
rect -4353 -1247 -4161 -1241
rect -4353 -1281 -4341 -1247
rect -4173 -1281 -4161 -1247
rect -4353 -1287 -4161 -1281
rect -4095 -1247 -3903 -1241
rect -4095 -1281 -4083 -1247
rect -3915 -1281 -3903 -1247
rect -4095 -1287 -3903 -1281
rect -3837 -1247 -3645 -1241
rect -3837 -1281 -3825 -1247
rect -3657 -1281 -3645 -1247
rect -3837 -1287 -3645 -1281
rect -3579 -1247 -3387 -1241
rect -3579 -1281 -3567 -1247
rect -3399 -1281 -3387 -1247
rect -3579 -1287 -3387 -1281
rect -3321 -1247 -3129 -1241
rect -3321 -1281 -3309 -1247
rect -3141 -1281 -3129 -1247
rect -3321 -1287 -3129 -1281
rect -3063 -1247 -2871 -1241
rect -3063 -1281 -3051 -1247
rect -2883 -1281 -2871 -1247
rect -3063 -1287 -2871 -1281
rect -2805 -1247 -2613 -1241
rect -2805 -1281 -2793 -1247
rect -2625 -1281 -2613 -1247
rect -2805 -1287 -2613 -1281
rect -2547 -1247 -2355 -1241
rect -2547 -1281 -2535 -1247
rect -2367 -1281 -2355 -1247
rect -2547 -1287 -2355 -1281
rect -2289 -1247 -2097 -1241
rect -2289 -1281 -2277 -1247
rect -2109 -1281 -2097 -1247
rect -2289 -1287 -2097 -1281
rect -2031 -1247 -1839 -1241
rect -2031 -1281 -2019 -1247
rect -1851 -1281 -1839 -1247
rect -2031 -1287 -1839 -1281
rect -1773 -1247 -1581 -1241
rect -1773 -1281 -1761 -1247
rect -1593 -1281 -1581 -1247
rect -1773 -1287 -1581 -1281
rect -1515 -1247 -1323 -1241
rect -1515 -1281 -1503 -1247
rect -1335 -1281 -1323 -1247
rect -1515 -1287 -1323 -1281
rect -1257 -1247 -1065 -1241
rect -1257 -1281 -1245 -1247
rect -1077 -1281 -1065 -1247
rect -1257 -1287 -1065 -1281
rect -999 -1247 -807 -1241
rect -999 -1281 -987 -1247
rect -819 -1281 -807 -1247
rect -999 -1287 -807 -1281
rect -741 -1247 -549 -1241
rect -741 -1281 -729 -1247
rect -561 -1281 -549 -1247
rect -741 -1287 -549 -1281
rect -483 -1247 -291 -1241
rect -483 -1281 -471 -1247
rect -303 -1281 -291 -1247
rect -483 -1287 -291 -1281
rect -225 -1247 -33 -1241
rect -225 -1281 -213 -1247
rect -45 -1281 -33 -1247
rect -225 -1287 -33 -1281
rect 33 -1247 225 -1241
rect 33 -1281 45 -1247
rect 213 -1281 225 -1247
rect 33 -1287 225 -1281
rect 291 -1247 483 -1241
rect 291 -1281 303 -1247
rect 471 -1281 483 -1247
rect 291 -1287 483 -1281
rect 549 -1247 741 -1241
rect 549 -1281 561 -1247
rect 729 -1281 741 -1247
rect 549 -1287 741 -1281
rect 807 -1247 999 -1241
rect 807 -1281 819 -1247
rect 987 -1281 999 -1247
rect 807 -1287 999 -1281
rect 1065 -1247 1257 -1241
rect 1065 -1281 1077 -1247
rect 1245 -1281 1257 -1247
rect 1065 -1287 1257 -1281
rect 1323 -1247 1515 -1241
rect 1323 -1281 1335 -1247
rect 1503 -1281 1515 -1247
rect 1323 -1287 1515 -1281
rect 1581 -1247 1773 -1241
rect 1581 -1281 1593 -1247
rect 1761 -1281 1773 -1247
rect 1581 -1287 1773 -1281
rect 1839 -1247 2031 -1241
rect 1839 -1281 1851 -1247
rect 2019 -1281 2031 -1247
rect 1839 -1287 2031 -1281
rect 2097 -1247 2289 -1241
rect 2097 -1281 2109 -1247
rect 2277 -1281 2289 -1247
rect 2097 -1287 2289 -1281
rect 2355 -1247 2547 -1241
rect 2355 -1281 2367 -1247
rect 2535 -1281 2547 -1247
rect 2355 -1287 2547 -1281
rect 2613 -1247 2805 -1241
rect 2613 -1281 2625 -1247
rect 2793 -1281 2805 -1247
rect 2613 -1287 2805 -1281
rect 2871 -1247 3063 -1241
rect 2871 -1281 2883 -1247
rect 3051 -1281 3063 -1247
rect 2871 -1287 3063 -1281
rect 3129 -1247 3321 -1241
rect 3129 -1281 3141 -1247
rect 3309 -1281 3321 -1247
rect 3129 -1287 3321 -1281
rect 3387 -1247 3579 -1241
rect 3387 -1281 3399 -1247
rect 3567 -1281 3579 -1247
rect 3387 -1287 3579 -1281
rect 3645 -1247 3837 -1241
rect 3645 -1281 3657 -1247
rect 3825 -1281 3837 -1247
rect 3645 -1287 3837 -1281
rect 3903 -1247 4095 -1241
rect 3903 -1281 3915 -1247
rect 4083 -1281 4095 -1247
rect 3903 -1287 4095 -1281
rect 4161 -1247 4353 -1241
rect 4161 -1281 4173 -1247
rect 4341 -1281 4353 -1247
rect 4161 -1287 4353 -1281
rect 4419 -1247 4611 -1241
rect 4419 -1281 4431 -1247
rect 4599 -1281 4611 -1247
rect 4419 -1287 4611 -1281
rect 4677 -1247 4869 -1241
rect 4677 -1281 4689 -1247
rect 4857 -1281 4869 -1247
rect 4677 -1287 4869 -1281
<< properties >>
string FIXED_BBOX -5036 -1402 5036 1402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 12 l 1 m 1 nf 38 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

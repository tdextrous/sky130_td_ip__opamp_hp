magic
tech sky130A
magscale 1 2
timestamp 1713300479
<< pwell >>
rect -2521 -1058 2521 1058
<< mvnmos >>
rect -2293 -800 -2093 800
rect -2035 -800 -1835 800
rect -1777 -800 -1577 800
rect -1519 -800 -1319 800
rect -1261 -800 -1061 800
rect -1003 -800 -803 800
rect -745 -800 -545 800
rect -487 -800 -287 800
rect -229 -800 -29 800
rect 29 -800 229 800
rect 287 -800 487 800
rect 545 -800 745 800
rect 803 -800 1003 800
rect 1061 -800 1261 800
rect 1319 -800 1519 800
rect 1577 -800 1777 800
rect 1835 -800 2035 800
rect 2093 -800 2293 800
<< mvndiff >>
rect -2351 788 -2293 800
rect -2351 -788 -2339 788
rect -2305 -788 -2293 788
rect -2351 -800 -2293 -788
rect -2093 788 -2035 800
rect -2093 -788 -2081 788
rect -2047 -788 -2035 788
rect -2093 -800 -2035 -788
rect -1835 788 -1777 800
rect -1835 -788 -1823 788
rect -1789 -788 -1777 788
rect -1835 -800 -1777 -788
rect -1577 788 -1519 800
rect -1577 -788 -1565 788
rect -1531 -788 -1519 788
rect -1577 -800 -1519 -788
rect -1319 788 -1261 800
rect -1319 -788 -1307 788
rect -1273 -788 -1261 788
rect -1319 -800 -1261 -788
rect -1061 788 -1003 800
rect -1061 -788 -1049 788
rect -1015 -788 -1003 788
rect -1061 -800 -1003 -788
rect -803 788 -745 800
rect -803 -788 -791 788
rect -757 -788 -745 788
rect -803 -800 -745 -788
rect -545 788 -487 800
rect -545 -788 -533 788
rect -499 -788 -487 788
rect -545 -800 -487 -788
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
rect 487 788 545 800
rect 487 -788 499 788
rect 533 -788 545 788
rect 487 -800 545 -788
rect 745 788 803 800
rect 745 -788 757 788
rect 791 -788 803 788
rect 745 -800 803 -788
rect 1003 788 1061 800
rect 1003 -788 1015 788
rect 1049 -788 1061 788
rect 1003 -800 1061 -788
rect 1261 788 1319 800
rect 1261 -788 1273 788
rect 1307 -788 1319 788
rect 1261 -800 1319 -788
rect 1519 788 1577 800
rect 1519 -788 1531 788
rect 1565 -788 1577 788
rect 1519 -800 1577 -788
rect 1777 788 1835 800
rect 1777 -788 1789 788
rect 1823 -788 1835 788
rect 1777 -800 1835 -788
rect 2035 788 2093 800
rect 2035 -788 2047 788
rect 2081 -788 2093 788
rect 2035 -800 2093 -788
rect 2293 788 2351 800
rect 2293 -788 2305 788
rect 2339 -788 2351 788
rect 2293 -800 2351 -788
<< mvndiffc >>
rect -2339 -788 -2305 788
rect -2081 -788 -2047 788
rect -1823 -788 -1789 788
rect -1565 -788 -1531 788
rect -1307 -788 -1273 788
rect -1049 -788 -1015 788
rect -791 -788 -757 788
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
rect 757 -788 791 788
rect 1015 -788 1049 788
rect 1273 -788 1307 788
rect 1531 -788 1565 788
rect 1789 -788 1823 788
rect 2047 -788 2081 788
rect 2305 -788 2339 788
<< mvpsubdiff >>
rect -2485 1010 2485 1022
rect -2485 976 -2377 1010
rect 2377 976 2485 1010
rect -2485 964 2485 976
rect -2485 914 -2427 964
rect -2485 -914 -2473 914
rect -2439 -914 -2427 914
rect 2427 914 2485 964
rect -2485 -964 -2427 -914
rect 2427 -914 2439 914
rect 2473 -914 2485 914
rect 2427 -964 2485 -914
rect -2485 -976 2485 -964
rect -2485 -1010 -2377 -976
rect 2377 -1010 2485 -976
rect -2485 -1022 2485 -1010
<< mvpsubdiffcont >>
rect -2377 976 2377 1010
rect -2473 -914 -2439 914
rect 2439 -914 2473 914
rect -2377 -1010 2377 -976
<< poly >>
rect -2259 872 -2127 888
rect -2259 855 -2243 872
rect -2293 838 -2243 855
rect -2143 855 -2127 872
rect -2001 872 -1869 888
rect -2001 855 -1985 872
rect -2143 838 -2093 855
rect -2293 800 -2093 838
rect -2035 838 -1985 855
rect -1885 855 -1869 872
rect -1743 872 -1611 888
rect -1743 855 -1727 872
rect -1885 838 -1835 855
rect -2035 800 -1835 838
rect -1777 838 -1727 855
rect -1627 855 -1611 872
rect -1485 872 -1353 888
rect -1485 855 -1469 872
rect -1627 838 -1577 855
rect -1777 800 -1577 838
rect -1519 838 -1469 855
rect -1369 855 -1353 872
rect -1227 872 -1095 888
rect -1227 855 -1211 872
rect -1369 838 -1319 855
rect -1519 800 -1319 838
rect -1261 838 -1211 855
rect -1111 855 -1095 872
rect -969 872 -837 888
rect -969 855 -953 872
rect -1111 838 -1061 855
rect -1261 800 -1061 838
rect -1003 838 -953 855
rect -853 855 -837 872
rect -711 872 -579 888
rect -711 855 -695 872
rect -853 838 -803 855
rect -1003 800 -803 838
rect -745 838 -695 855
rect -595 855 -579 872
rect -453 872 -321 888
rect -453 855 -437 872
rect -595 838 -545 855
rect -745 800 -545 838
rect -487 838 -437 855
rect -337 855 -321 872
rect -195 872 -63 888
rect -195 855 -179 872
rect -337 838 -287 855
rect -487 800 -287 838
rect -229 838 -179 855
rect -79 855 -63 872
rect 63 872 195 888
rect 63 855 79 872
rect -79 838 -29 855
rect -229 800 -29 838
rect 29 838 79 855
rect 179 855 195 872
rect 321 872 453 888
rect 321 855 337 872
rect 179 838 229 855
rect 29 800 229 838
rect 287 838 337 855
rect 437 855 453 872
rect 579 872 711 888
rect 579 855 595 872
rect 437 838 487 855
rect 287 800 487 838
rect 545 838 595 855
rect 695 855 711 872
rect 837 872 969 888
rect 837 855 853 872
rect 695 838 745 855
rect 545 800 745 838
rect 803 838 853 855
rect 953 855 969 872
rect 1095 872 1227 888
rect 1095 855 1111 872
rect 953 838 1003 855
rect 803 800 1003 838
rect 1061 838 1111 855
rect 1211 855 1227 872
rect 1353 872 1485 888
rect 1353 855 1369 872
rect 1211 838 1261 855
rect 1061 800 1261 838
rect 1319 838 1369 855
rect 1469 855 1485 872
rect 1611 872 1743 888
rect 1611 855 1627 872
rect 1469 838 1519 855
rect 1319 800 1519 838
rect 1577 838 1627 855
rect 1727 855 1743 872
rect 1869 872 2001 888
rect 1869 855 1885 872
rect 1727 838 1777 855
rect 1577 800 1777 838
rect 1835 838 1885 855
rect 1985 855 2001 872
rect 2127 872 2259 888
rect 2127 855 2143 872
rect 1985 838 2035 855
rect 1835 800 2035 838
rect 2093 838 2143 855
rect 2243 855 2259 872
rect 2243 838 2293 855
rect 2093 800 2293 838
rect -2293 -838 -2093 -800
rect -2293 -855 -2243 -838
rect -2259 -872 -2243 -855
rect -2143 -855 -2093 -838
rect -2035 -838 -1835 -800
rect -2035 -855 -1985 -838
rect -2143 -872 -2127 -855
rect -2259 -888 -2127 -872
rect -2001 -872 -1985 -855
rect -1885 -855 -1835 -838
rect -1777 -838 -1577 -800
rect -1777 -855 -1727 -838
rect -1885 -872 -1869 -855
rect -2001 -888 -1869 -872
rect -1743 -872 -1727 -855
rect -1627 -855 -1577 -838
rect -1519 -838 -1319 -800
rect -1519 -855 -1469 -838
rect -1627 -872 -1611 -855
rect -1743 -888 -1611 -872
rect -1485 -872 -1469 -855
rect -1369 -855 -1319 -838
rect -1261 -838 -1061 -800
rect -1261 -855 -1211 -838
rect -1369 -872 -1353 -855
rect -1485 -888 -1353 -872
rect -1227 -872 -1211 -855
rect -1111 -855 -1061 -838
rect -1003 -838 -803 -800
rect -1003 -855 -953 -838
rect -1111 -872 -1095 -855
rect -1227 -888 -1095 -872
rect -969 -872 -953 -855
rect -853 -855 -803 -838
rect -745 -838 -545 -800
rect -745 -855 -695 -838
rect -853 -872 -837 -855
rect -969 -888 -837 -872
rect -711 -872 -695 -855
rect -595 -855 -545 -838
rect -487 -838 -287 -800
rect -487 -855 -437 -838
rect -595 -872 -579 -855
rect -711 -888 -579 -872
rect -453 -872 -437 -855
rect -337 -855 -287 -838
rect -229 -838 -29 -800
rect -229 -855 -179 -838
rect -337 -872 -321 -855
rect -453 -888 -321 -872
rect -195 -872 -179 -855
rect -79 -855 -29 -838
rect 29 -838 229 -800
rect 29 -855 79 -838
rect -79 -872 -63 -855
rect -195 -888 -63 -872
rect 63 -872 79 -855
rect 179 -855 229 -838
rect 287 -838 487 -800
rect 287 -855 337 -838
rect 179 -872 195 -855
rect 63 -888 195 -872
rect 321 -872 337 -855
rect 437 -855 487 -838
rect 545 -838 745 -800
rect 545 -855 595 -838
rect 437 -872 453 -855
rect 321 -888 453 -872
rect 579 -872 595 -855
rect 695 -855 745 -838
rect 803 -838 1003 -800
rect 803 -855 853 -838
rect 695 -872 711 -855
rect 579 -888 711 -872
rect 837 -872 853 -855
rect 953 -855 1003 -838
rect 1061 -838 1261 -800
rect 1061 -855 1111 -838
rect 953 -872 969 -855
rect 837 -888 969 -872
rect 1095 -872 1111 -855
rect 1211 -855 1261 -838
rect 1319 -838 1519 -800
rect 1319 -855 1369 -838
rect 1211 -872 1227 -855
rect 1095 -888 1227 -872
rect 1353 -872 1369 -855
rect 1469 -855 1519 -838
rect 1577 -838 1777 -800
rect 1577 -855 1627 -838
rect 1469 -872 1485 -855
rect 1353 -888 1485 -872
rect 1611 -872 1627 -855
rect 1727 -855 1777 -838
rect 1835 -838 2035 -800
rect 1835 -855 1885 -838
rect 1727 -872 1743 -855
rect 1611 -888 1743 -872
rect 1869 -872 1885 -855
rect 1985 -855 2035 -838
rect 2093 -838 2293 -800
rect 2093 -855 2143 -838
rect 1985 -872 2001 -855
rect 1869 -888 2001 -872
rect 2127 -872 2143 -855
rect 2243 -855 2293 -838
rect 2243 -872 2259 -855
rect 2127 -888 2259 -872
<< polycont >>
rect -2243 838 -2143 872
rect -1985 838 -1885 872
rect -1727 838 -1627 872
rect -1469 838 -1369 872
rect -1211 838 -1111 872
rect -953 838 -853 872
rect -695 838 -595 872
rect -437 838 -337 872
rect -179 838 -79 872
rect 79 838 179 872
rect 337 838 437 872
rect 595 838 695 872
rect 853 838 953 872
rect 1111 838 1211 872
rect 1369 838 1469 872
rect 1627 838 1727 872
rect 1885 838 1985 872
rect 2143 838 2243 872
rect -2243 -872 -2143 -838
rect -1985 -872 -1885 -838
rect -1727 -872 -1627 -838
rect -1469 -872 -1369 -838
rect -1211 -872 -1111 -838
rect -953 -872 -853 -838
rect -695 -872 -595 -838
rect -437 -872 -337 -838
rect -179 -872 -79 -838
rect 79 -872 179 -838
rect 337 -872 437 -838
rect 595 -872 695 -838
rect 853 -872 953 -838
rect 1111 -872 1211 -838
rect 1369 -872 1469 -838
rect 1627 -872 1727 -838
rect 1885 -872 1985 -838
rect 2143 -872 2243 -838
<< locali >>
rect -2473 976 -2377 1010
rect 2377 976 2473 1010
rect -2473 914 -2439 976
rect 2439 914 2473 976
rect -2259 838 -2243 872
rect -2143 838 -2127 872
rect -2001 838 -1985 872
rect -1885 838 -1869 872
rect -1743 838 -1727 872
rect -1627 838 -1611 872
rect -1485 838 -1469 872
rect -1369 838 -1353 872
rect -1227 838 -1211 872
rect -1111 838 -1095 872
rect -969 838 -953 872
rect -853 838 -837 872
rect -711 838 -695 872
rect -595 838 -579 872
rect -453 838 -437 872
rect -337 838 -321 872
rect -195 838 -179 872
rect -79 838 -63 872
rect 63 838 79 872
rect 179 838 195 872
rect 321 838 337 872
rect 437 838 453 872
rect 579 838 595 872
rect 695 838 711 872
rect 837 838 853 872
rect 953 838 969 872
rect 1095 838 1111 872
rect 1211 838 1227 872
rect 1353 838 1369 872
rect 1469 838 1485 872
rect 1611 838 1627 872
rect 1727 838 1743 872
rect 1869 838 1885 872
rect 1985 838 2001 872
rect 2127 838 2143 872
rect 2243 838 2259 872
rect -2339 788 -2305 804
rect -2339 -804 -2305 -788
rect -2081 788 -2047 804
rect -2081 -804 -2047 -788
rect -1823 788 -1789 804
rect -1823 -804 -1789 -788
rect -1565 788 -1531 804
rect -1565 -804 -1531 -788
rect -1307 788 -1273 804
rect -1307 -804 -1273 -788
rect -1049 788 -1015 804
rect -1049 -804 -1015 -788
rect -791 788 -757 804
rect -791 -804 -757 -788
rect -533 788 -499 804
rect -533 -804 -499 -788
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
rect 499 788 533 804
rect 499 -804 533 -788
rect 757 788 791 804
rect 757 -804 791 -788
rect 1015 788 1049 804
rect 1015 -804 1049 -788
rect 1273 788 1307 804
rect 1273 -804 1307 -788
rect 1531 788 1565 804
rect 1531 -804 1565 -788
rect 1789 788 1823 804
rect 1789 -804 1823 -788
rect 2047 788 2081 804
rect 2047 -804 2081 -788
rect 2305 788 2339 804
rect 2305 -804 2339 -788
rect -2259 -872 -2243 -838
rect -2143 -872 -2127 -838
rect -2001 -872 -1985 -838
rect -1885 -872 -1869 -838
rect -1743 -872 -1727 -838
rect -1627 -872 -1611 -838
rect -1485 -872 -1469 -838
rect -1369 -872 -1353 -838
rect -1227 -872 -1211 -838
rect -1111 -872 -1095 -838
rect -969 -872 -953 -838
rect -853 -872 -837 -838
rect -711 -872 -695 -838
rect -595 -872 -579 -838
rect -453 -872 -437 -838
rect -337 -872 -321 -838
rect -195 -872 -179 -838
rect -79 -872 -63 -838
rect 63 -872 79 -838
rect 179 -872 195 -838
rect 321 -872 337 -838
rect 437 -872 453 -838
rect 579 -872 595 -838
rect 695 -872 711 -838
rect 837 -872 853 -838
rect 953 -872 969 -838
rect 1095 -872 1111 -838
rect 1211 -872 1227 -838
rect 1353 -872 1369 -838
rect 1469 -872 1485 -838
rect 1611 -872 1627 -838
rect 1727 -872 1743 -838
rect 1869 -872 1885 -838
rect 1985 -872 2001 -838
rect 2127 -872 2143 -838
rect 2243 -872 2259 -838
rect -2473 -976 -2439 -914
rect 2439 -976 2473 -914
rect -2473 -1010 -2377 -976
rect 2377 -1010 2473 -976
<< viali >>
rect -2243 838 -2143 872
rect -1985 838 -1885 872
rect -1727 838 -1627 872
rect -1469 838 -1369 872
rect -1211 838 -1111 872
rect -953 838 -853 872
rect -695 838 -595 872
rect -437 838 -337 872
rect -179 838 -79 872
rect 79 838 179 872
rect 337 838 437 872
rect 595 838 695 872
rect 853 838 953 872
rect 1111 838 1211 872
rect 1369 838 1469 872
rect 1627 838 1727 872
rect 1885 838 1985 872
rect 2143 838 2243 872
rect -2339 -788 -2305 788
rect -2081 -788 -2047 788
rect -1823 -788 -1789 788
rect -1565 -788 -1531 788
rect -1307 -788 -1273 788
rect -1049 -788 -1015 788
rect -791 -788 -757 788
rect -533 -788 -499 788
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
rect 499 -788 533 788
rect 757 -788 791 788
rect 1015 -788 1049 788
rect 1273 -788 1307 788
rect 1531 -788 1565 788
rect 1789 -788 1823 788
rect 2047 -788 2081 788
rect 2305 -788 2339 788
rect -2243 -872 -2143 -838
rect -1985 -872 -1885 -838
rect -1727 -872 -1627 -838
rect -1469 -872 -1369 -838
rect -1211 -872 -1111 -838
rect -953 -872 -853 -838
rect -695 -872 -595 -838
rect -437 -872 -337 -838
rect -179 -872 -79 -838
rect 79 -872 179 -838
rect 337 -872 437 -838
rect 595 -872 695 -838
rect 853 -872 953 -838
rect 1111 -872 1211 -838
rect 1369 -872 1469 -838
rect 1627 -872 1727 -838
rect 1885 -872 1985 -838
rect 2143 -872 2243 -838
<< metal1 >>
rect -2255 872 -2131 878
rect -2255 838 -2243 872
rect -2143 838 -2131 872
rect -2255 832 -2131 838
rect -1997 872 -1873 878
rect -1997 838 -1985 872
rect -1885 838 -1873 872
rect -1997 832 -1873 838
rect -1739 872 -1615 878
rect -1739 838 -1727 872
rect -1627 838 -1615 872
rect -1739 832 -1615 838
rect -1481 872 -1357 878
rect -1481 838 -1469 872
rect -1369 838 -1357 872
rect -1481 832 -1357 838
rect -1223 872 -1099 878
rect -1223 838 -1211 872
rect -1111 838 -1099 872
rect -1223 832 -1099 838
rect -965 872 -841 878
rect -965 838 -953 872
rect -853 838 -841 872
rect -965 832 -841 838
rect -707 872 -583 878
rect -707 838 -695 872
rect -595 838 -583 872
rect -707 832 -583 838
rect -449 872 -325 878
rect -449 838 -437 872
rect -337 838 -325 872
rect -449 832 -325 838
rect -191 872 -67 878
rect -191 838 -179 872
rect -79 838 -67 872
rect -191 832 -67 838
rect 67 872 191 878
rect 67 838 79 872
rect 179 838 191 872
rect 67 832 191 838
rect 325 872 449 878
rect 325 838 337 872
rect 437 838 449 872
rect 325 832 449 838
rect 583 872 707 878
rect 583 838 595 872
rect 695 838 707 872
rect 583 832 707 838
rect 841 872 965 878
rect 841 838 853 872
rect 953 838 965 872
rect 841 832 965 838
rect 1099 872 1223 878
rect 1099 838 1111 872
rect 1211 838 1223 872
rect 1099 832 1223 838
rect 1357 872 1481 878
rect 1357 838 1369 872
rect 1469 838 1481 872
rect 1357 832 1481 838
rect 1615 872 1739 878
rect 1615 838 1627 872
rect 1727 838 1739 872
rect 1615 832 1739 838
rect 1873 872 1997 878
rect 1873 838 1885 872
rect 1985 838 1997 872
rect 1873 832 1997 838
rect 2131 872 2255 878
rect 2131 838 2143 872
rect 2243 838 2255 872
rect 2131 832 2255 838
rect -2345 788 -2299 800
rect -2345 -788 -2339 788
rect -2305 -788 -2299 788
rect -2345 -800 -2299 -788
rect -2087 788 -2041 800
rect -2087 -788 -2081 788
rect -2047 -788 -2041 788
rect -2087 -800 -2041 -788
rect -1829 788 -1783 800
rect -1829 -788 -1823 788
rect -1789 -788 -1783 788
rect -1829 -800 -1783 -788
rect -1571 788 -1525 800
rect -1571 -788 -1565 788
rect -1531 -788 -1525 788
rect -1571 -800 -1525 -788
rect -1313 788 -1267 800
rect -1313 -788 -1307 788
rect -1273 -788 -1267 788
rect -1313 -800 -1267 -788
rect -1055 788 -1009 800
rect -1055 -788 -1049 788
rect -1015 -788 -1009 788
rect -1055 -800 -1009 -788
rect -797 788 -751 800
rect -797 -788 -791 788
rect -757 -788 -751 788
rect -797 -800 -751 -788
rect -539 788 -493 800
rect -539 -788 -533 788
rect -499 -788 -493 788
rect -539 -800 -493 -788
rect -281 788 -235 800
rect -281 -788 -275 788
rect -241 -788 -235 788
rect -281 -800 -235 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 235 788 281 800
rect 235 -788 241 788
rect 275 -788 281 788
rect 235 -800 281 -788
rect 493 788 539 800
rect 493 -788 499 788
rect 533 -788 539 788
rect 493 -800 539 -788
rect 751 788 797 800
rect 751 -788 757 788
rect 791 -788 797 788
rect 751 -800 797 -788
rect 1009 788 1055 800
rect 1009 -788 1015 788
rect 1049 -788 1055 788
rect 1009 -800 1055 -788
rect 1267 788 1313 800
rect 1267 -788 1273 788
rect 1307 -788 1313 788
rect 1267 -800 1313 -788
rect 1525 788 1571 800
rect 1525 -788 1531 788
rect 1565 -788 1571 788
rect 1525 -800 1571 -788
rect 1783 788 1829 800
rect 1783 -788 1789 788
rect 1823 -788 1829 788
rect 1783 -800 1829 -788
rect 2041 788 2087 800
rect 2041 -788 2047 788
rect 2081 -788 2087 788
rect 2041 -800 2087 -788
rect 2299 788 2345 800
rect 2299 -788 2305 788
rect 2339 -788 2345 788
rect 2299 -800 2345 -788
rect -2255 -838 -2131 -832
rect -2255 -872 -2243 -838
rect -2143 -872 -2131 -838
rect -2255 -878 -2131 -872
rect -1997 -838 -1873 -832
rect -1997 -872 -1985 -838
rect -1885 -872 -1873 -838
rect -1997 -878 -1873 -872
rect -1739 -838 -1615 -832
rect -1739 -872 -1727 -838
rect -1627 -872 -1615 -838
rect -1739 -878 -1615 -872
rect -1481 -838 -1357 -832
rect -1481 -872 -1469 -838
rect -1369 -872 -1357 -838
rect -1481 -878 -1357 -872
rect -1223 -838 -1099 -832
rect -1223 -872 -1211 -838
rect -1111 -872 -1099 -838
rect -1223 -878 -1099 -872
rect -965 -838 -841 -832
rect -965 -872 -953 -838
rect -853 -872 -841 -838
rect -965 -878 -841 -872
rect -707 -838 -583 -832
rect -707 -872 -695 -838
rect -595 -872 -583 -838
rect -707 -878 -583 -872
rect -449 -838 -325 -832
rect -449 -872 -437 -838
rect -337 -872 -325 -838
rect -449 -878 -325 -872
rect -191 -838 -67 -832
rect -191 -872 -179 -838
rect -79 -872 -67 -838
rect -191 -878 -67 -872
rect 67 -838 191 -832
rect 67 -872 79 -838
rect 179 -872 191 -838
rect 67 -878 191 -872
rect 325 -838 449 -832
rect 325 -872 337 -838
rect 437 -872 449 -838
rect 325 -878 449 -872
rect 583 -838 707 -832
rect 583 -872 595 -838
rect 695 -872 707 -838
rect 583 -878 707 -872
rect 841 -838 965 -832
rect 841 -872 853 -838
rect 953 -872 965 -838
rect 841 -878 965 -872
rect 1099 -838 1223 -832
rect 1099 -872 1111 -838
rect 1211 -872 1223 -838
rect 1099 -878 1223 -872
rect 1357 -838 1481 -832
rect 1357 -872 1369 -838
rect 1469 -872 1481 -838
rect 1357 -878 1481 -872
rect 1615 -838 1739 -832
rect 1615 -872 1627 -838
rect 1727 -872 1739 -838
rect 1615 -878 1739 -872
rect 1873 -838 1997 -832
rect 1873 -872 1885 -838
rect 1985 -872 1997 -838
rect 1873 -878 1997 -872
rect 2131 -838 2255 -832
rect 2131 -872 2143 -838
rect 2243 -872 2255 -838
rect 2131 -878 2255 -872
<< properties >>
string FIXED_BBOX -2456 -993 2456 993
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 1 m 1 nf 18 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

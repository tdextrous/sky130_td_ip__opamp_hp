magic
tech sky130A
magscale 1 2
timestamp 1713416651
<< error_p >>
rect -743 481 -679 487
rect -585 481 -521 487
rect -427 481 -363 487
rect -269 481 -205 487
rect -111 481 -47 487
rect 47 481 111 487
rect 205 481 269 487
rect 363 481 427 487
rect 521 481 585 487
rect 679 481 743 487
rect -743 447 -731 481
rect -585 447 -573 481
rect -427 447 -415 481
rect -269 447 -257 481
rect -111 447 -99 481
rect 47 447 59 481
rect 205 447 217 481
rect 363 447 375 481
rect 521 447 533 481
rect 679 447 691 481
rect -743 441 -679 447
rect -585 441 -521 447
rect -427 441 -363 447
rect -269 441 -205 447
rect -111 441 -47 447
rect 47 441 111 447
rect 205 441 269 447
rect 363 441 427 447
rect 521 441 585 447
rect 679 441 743 447
rect -743 -447 -679 -441
rect -585 -447 -521 -441
rect -427 -447 -363 -441
rect -269 -447 -205 -441
rect -111 -447 -47 -441
rect 47 -447 111 -441
rect 205 -447 269 -441
rect 363 -447 427 -441
rect 521 -447 585 -441
rect 679 -447 743 -441
rect -743 -481 -731 -447
rect -585 -481 -573 -447
rect -427 -481 -415 -447
rect -269 -481 -257 -447
rect -111 -481 -99 -447
rect 47 -481 59 -447
rect 205 -481 217 -447
rect 363 -481 375 -447
rect 521 -481 533 -447
rect 679 -481 691 -447
rect -743 -487 -679 -481
rect -585 -487 -521 -481
rect -427 -487 -363 -481
rect -269 -487 -205 -481
rect -111 -487 -47 -481
rect 47 -487 111 -481
rect 205 -487 269 -481
rect 363 -487 427 -481
rect 521 -487 585 -481
rect 679 -487 743 -481
<< nwell >>
rect -1019 -697 1019 697
<< mvpmos >>
rect -761 -400 -661 400
rect -603 -400 -503 400
rect -445 -400 -345 400
rect -287 -400 -187 400
rect -129 -400 -29 400
rect 29 -400 129 400
rect 187 -400 287 400
rect 345 -400 445 400
rect 503 -400 603 400
rect 661 -400 761 400
<< mvpdiff >>
rect -819 388 -761 400
rect -819 -388 -807 388
rect -773 -388 -761 388
rect -819 -400 -761 -388
rect -661 388 -603 400
rect -661 -388 -649 388
rect -615 -388 -603 388
rect -661 -400 -603 -388
rect -503 388 -445 400
rect -503 -388 -491 388
rect -457 -388 -445 388
rect -503 -400 -445 -388
rect -345 388 -287 400
rect -345 -388 -333 388
rect -299 -388 -287 388
rect -345 -400 -287 -388
rect -187 388 -129 400
rect -187 -388 -175 388
rect -141 -388 -129 388
rect -187 -400 -129 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 129 388 187 400
rect 129 -388 141 388
rect 175 -388 187 388
rect 129 -400 187 -388
rect 287 388 345 400
rect 287 -388 299 388
rect 333 -388 345 388
rect 287 -400 345 -388
rect 445 388 503 400
rect 445 -388 457 388
rect 491 -388 503 388
rect 445 -400 503 -388
rect 603 388 661 400
rect 603 -388 615 388
rect 649 -388 661 388
rect 603 -400 661 -388
rect 761 388 819 400
rect 761 -388 773 388
rect 807 -388 819 388
rect 761 -400 819 -388
<< mvpdiffc >>
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
<< mvnsubdiff >>
rect -953 619 953 631
rect -953 585 -845 619
rect 845 585 953 619
rect -953 573 953 585
rect -953 523 -895 573
rect -953 -523 -941 523
rect -907 -523 -895 523
rect 895 523 953 573
rect -953 -573 -895 -523
rect 895 -523 907 523
rect 941 -523 953 523
rect 895 -573 953 -523
rect -953 -585 953 -573
rect -953 -619 -845 -585
rect 845 -619 953 -585
rect -953 -631 953 -619
<< mvnsubdiffcont >>
rect -845 585 845 619
rect -941 -523 -907 523
rect 907 -523 941 523
rect -845 -619 845 -585
<< poly >>
rect -747 481 -675 497
rect -747 464 -731 481
rect -761 447 -731 464
rect -691 464 -675 481
rect -589 481 -517 497
rect -589 464 -573 481
rect -691 447 -661 464
rect -761 400 -661 447
rect -603 447 -573 464
rect -533 464 -517 481
rect -431 481 -359 497
rect -431 464 -415 481
rect -533 447 -503 464
rect -603 400 -503 447
rect -445 447 -415 464
rect -375 464 -359 481
rect -273 481 -201 497
rect -273 464 -257 481
rect -375 447 -345 464
rect -445 400 -345 447
rect -287 447 -257 464
rect -217 464 -201 481
rect -115 481 -43 497
rect -115 464 -99 481
rect -217 447 -187 464
rect -287 400 -187 447
rect -129 447 -99 464
rect -59 464 -43 481
rect 43 481 115 497
rect 43 464 59 481
rect -59 447 -29 464
rect -129 400 -29 447
rect 29 447 59 464
rect 99 464 115 481
rect 201 481 273 497
rect 201 464 217 481
rect 99 447 129 464
rect 29 400 129 447
rect 187 447 217 464
rect 257 464 273 481
rect 359 481 431 497
rect 359 464 375 481
rect 257 447 287 464
rect 187 400 287 447
rect 345 447 375 464
rect 415 464 431 481
rect 517 481 589 497
rect 517 464 533 481
rect 415 447 445 464
rect 345 400 445 447
rect 503 447 533 464
rect 573 464 589 481
rect 675 481 747 497
rect 675 464 691 481
rect 573 447 603 464
rect 503 400 603 447
rect 661 447 691 464
rect 731 464 747 481
rect 731 447 761 464
rect 661 400 761 447
rect -761 -447 -661 -400
rect -761 -464 -731 -447
rect -747 -481 -731 -464
rect -691 -464 -661 -447
rect -603 -447 -503 -400
rect -603 -464 -573 -447
rect -691 -481 -675 -464
rect -747 -497 -675 -481
rect -589 -481 -573 -464
rect -533 -464 -503 -447
rect -445 -447 -345 -400
rect -445 -464 -415 -447
rect -533 -481 -517 -464
rect -589 -497 -517 -481
rect -431 -481 -415 -464
rect -375 -464 -345 -447
rect -287 -447 -187 -400
rect -287 -464 -257 -447
rect -375 -481 -359 -464
rect -431 -497 -359 -481
rect -273 -481 -257 -464
rect -217 -464 -187 -447
rect -129 -447 -29 -400
rect -129 -464 -99 -447
rect -217 -481 -201 -464
rect -273 -497 -201 -481
rect -115 -481 -99 -464
rect -59 -464 -29 -447
rect 29 -447 129 -400
rect 29 -464 59 -447
rect -59 -481 -43 -464
rect -115 -497 -43 -481
rect 43 -481 59 -464
rect 99 -464 129 -447
rect 187 -447 287 -400
rect 187 -464 217 -447
rect 99 -481 115 -464
rect 43 -497 115 -481
rect 201 -481 217 -464
rect 257 -464 287 -447
rect 345 -447 445 -400
rect 345 -464 375 -447
rect 257 -481 273 -464
rect 201 -497 273 -481
rect 359 -481 375 -464
rect 415 -464 445 -447
rect 503 -447 603 -400
rect 503 -464 533 -447
rect 415 -481 431 -464
rect 359 -497 431 -481
rect 517 -481 533 -464
rect 573 -464 603 -447
rect 661 -447 761 -400
rect 661 -464 691 -447
rect 573 -481 589 -464
rect 517 -497 589 -481
rect 675 -481 691 -464
rect 731 -464 761 -447
rect 731 -481 747 -464
rect 675 -497 747 -481
<< polycont >>
rect -731 447 -691 481
rect -573 447 -533 481
rect -415 447 -375 481
rect -257 447 -217 481
rect -99 447 -59 481
rect 59 447 99 481
rect 217 447 257 481
rect 375 447 415 481
rect 533 447 573 481
rect 691 447 731 481
rect -731 -481 -691 -447
rect -573 -481 -533 -447
rect -415 -481 -375 -447
rect -257 -481 -217 -447
rect -99 -481 -59 -447
rect 59 -481 99 -447
rect 217 -481 257 -447
rect 375 -481 415 -447
rect 533 -481 573 -447
rect 691 -481 731 -447
<< locali >>
rect -941 585 -845 619
rect 845 585 941 619
rect -941 523 -907 585
rect 907 523 941 585
rect -747 447 -731 481
rect -691 447 -675 481
rect -589 447 -573 481
rect -533 447 -517 481
rect -431 447 -415 481
rect -375 447 -359 481
rect -273 447 -257 481
rect -217 447 -201 481
rect -115 447 -99 481
rect -59 447 -43 481
rect 43 447 59 481
rect 99 447 115 481
rect 201 447 217 481
rect 257 447 273 481
rect 359 447 375 481
rect 415 447 431 481
rect 517 447 533 481
rect 573 447 589 481
rect 675 447 691 481
rect 731 447 747 481
rect -807 388 -773 404
rect -807 -404 -773 -388
rect -649 388 -615 404
rect -649 -404 -615 -388
rect -491 388 -457 404
rect -491 -404 -457 -388
rect -333 388 -299 404
rect -333 -404 -299 -388
rect -175 388 -141 404
rect -175 -404 -141 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 141 388 175 404
rect 141 -404 175 -388
rect 299 388 333 404
rect 299 -404 333 -388
rect 457 388 491 404
rect 457 -404 491 -388
rect 615 388 649 404
rect 615 -404 649 -388
rect 773 388 807 404
rect 773 -404 807 -388
rect -747 -481 -731 -447
rect -691 -481 -675 -447
rect -589 -481 -573 -447
rect -533 -481 -517 -447
rect -431 -481 -415 -447
rect -375 -481 -359 -447
rect -273 -481 -257 -447
rect -217 -481 -201 -447
rect -115 -481 -99 -447
rect -59 -481 -43 -447
rect 43 -481 59 -447
rect 99 -481 115 -447
rect 201 -481 217 -447
rect 257 -481 273 -447
rect 359 -481 375 -447
rect 415 -481 431 -447
rect 517 -481 533 -447
rect 573 -481 589 -447
rect 675 -481 691 -447
rect 731 -481 747 -447
rect -941 -585 -907 -523
rect 907 -585 941 -523
rect -941 -619 -845 -585
rect 845 -619 941 -585
<< viali >>
rect -731 447 -691 481
rect -573 447 -533 481
rect -415 447 -375 481
rect -257 447 -217 481
rect -99 447 -59 481
rect 59 447 99 481
rect 217 447 257 481
rect 375 447 415 481
rect 533 447 573 481
rect 691 447 731 481
rect -807 -388 -773 388
rect -649 -388 -615 388
rect -491 -388 -457 388
rect -333 -388 -299 388
rect -175 -388 -141 388
rect -17 -388 17 388
rect 141 -388 175 388
rect 299 -388 333 388
rect 457 -388 491 388
rect 615 -388 649 388
rect 773 -388 807 388
rect -731 -481 -691 -447
rect -573 -481 -533 -447
rect -415 -481 -375 -447
rect -257 -481 -217 -447
rect -99 -481 -59 -447
rect 59 -481 99 -447
rect 217 -481 257 -447
rect 375 -481 415 -447
rect 533 -481 573 -447
rect 691 -481 731 -447
<< metal1 >>
rect -743 481 -679 487
rect -743 447 -731 481
rect -691 447 -679 481
rect -743 441 -679 447
rect -585 481 -521 487
rect -585 447 -573 481
rect -533 447 -521 481
rect -585 441 -521 447
rect -427 481 -363 487
rect -427 447 -415 481
rect -375 447 -363 481
rect -427 441 -363 447
rect -269 481 -205 487
rect -269 447 -257 481
rect -217 447 -205 481
rect -269 441 -205 447
rect -111 481 -47 487
rect -111 447 -99 481
rect -59 447 -47 481
rect -111 441 -47 447
rect 47 481 111 487
rect 47 447 59 481
rect 99 447 111 481
rect 47 441 111 447
rect 205 481 269 487
rect 205 447 217 481
rect 257 447 269 481
rect 205 441 269 447
rect 363 481 427 487
rect 363 447 375 481
rect 415 447 427 481
rect 363 441 427 447
rect 521 481 585 487
rect 521 447 533 481
rect 573 447 585 481
rect 521 441 585 447
rect 679 481 743 487
rect 679 447 691 481
rect 731 447 743 481
rect 679 441 743 447
rect -813 388 -767 400
rect -813 -388 -807 388
rect -773 -388 -767 388
rect -813 -400 -767 -388
rect -655 388 -609 400
rect -655 -388 -649 388
rect -615 -388 -609 388
rect -655 -400 -609 -388
rect -497 388 -451 400
rect -497 -388 -491 388
rect -457 -388 -451 388
rect -497 -400 -451 -388
rect -339 388 -293 400
rect -339 -388 -333 388
rect -299 -388 -293 388
rect -339 -400 -293 -388
rect -181 388 -135 400
rect -181 -388 -175 388
rect -141 -388 -135 388
rect -181 -400 -135 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 135 388 181 400
rect 135 -388 141 388
rect 175 -388 181 388
rect 135 -400 181 -388
rect 293 388 339 400
rect 293 -388 299 388
rect 333 -388 339 388
rect 293 -400 339 -388
rect 451 388 497 400
rect 451 -388 457 388
rect 491 -388 497 388
rect 451 -400 497 -388
rect 609 388 655 400
rect 609 -388 615 388
rect 649 -388 655 388
rect 609 -400 655 -388
rect 767 388 813 400
rect 767 -388 773 388
rect 807 -388 813 388
rect 767 -400 813 -388
rect -743 -447 -679 -441
rect -743 -481 -731 -447
rect -691 -481 -679 -447
rect -743 -487 -679 -481
rect -585 -447 -521 -441
rect -585 -481 -573 -447
rect -533 -481 -521 -447
rect -585 -487 -521 -481
rect -427 -447 -363 -441
rect -427 -481 -415 -447
rect -375 -481 -363 -447
rect -427 -487 -363 -481
rect -269 -447 -205 -441
rect -269 -481 -257 -447
rect -217 -481 -205 -447
rect -269 -487 -205 -481
rect -111 -447 -47 -441
rect -111 -481 -99 -447
rect -59 -481 -47 -447
rect -111 -487 -47 -481
rect 47 -447 111 -441
rect 47 -481 59 -447
rect 99 -481 111 -447
rect 47 -487 111 -481
rect 205 -447 269 -441
rect 205 -481 217 -447
rect 257 -481 269 -447
rect 205 -487 269 -481
rect 363 -447 427 -441
rect 363 -481 375 -447
rect 415 -481 427 -447
rect 363 -487 427 -481
rect 521 -447 585 -441
rect 521 -481 533 -447
rect 573 -481 585 -447
rect 521 -487 585 -481
rect 679 -447 743 -441
rect 679 -481 691 -447
rect 731 -481 743 -447
rect 679 -487 743 -481
<< properties >>
string FIXED_BBOX -924 -602 924 602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 0.5 m 1 nf 10 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

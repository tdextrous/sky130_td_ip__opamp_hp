magic
tech sky130A
magscale 1 2
timestamp 1713235147
<< metal3 >>
rect -15128 4492 -11556 4520
rect -15128 2468 -11640 4492
rect -11576 2468 -11556 4492
rect -15128 2440 -11556 2468
rect -11316 4492 -7744 4520
rect -11316 2468 -7828 4492
rect -7764 2468 -7744 4492
rect -11316 2440 -7744 2468
rect -7504 4492 -3932 4520
rect -7504 2468 -4016 4492
rect -3952 2468 -3932 4492
rect -7504 2440 -3932 2468
rect -3692 4492 -120 4520
rect -3692 2468 -204 4492
rect -140 2468 -120 4492
rect -3692 2440 -120 2468
rect 120 4492 3692 4520
rect 120 2468 3608 4492
rect 3672 2468 3692 4492
rect 120 2440 3692 2468
rect 3932 4492 7504 4520
rect 3932 2468 7420 4492
rect 7484 2468 7504 4492
rect 3932 2440 7504 2468
rect 7744 4492 11316 4520
rect 7744 2468 11232 4492
rect 11296 2468 11316 4492
rect 7744 2440 11316 2468
rect 11556 4492 15128 4520
rect 11556 2468 15044 4492
rect 15108 2468 15128 4492
rect 11556 2440 15128 2468
rect -15128 2172 -11556 2200
rect -15128 148 -11640 2172
rect -11576 148 -11556 2172
rect -15128 120 -11556 148
rect -11316 2172 -7744 2200
rect -11316 148 -7828 2172
rect -7764 148 -7744 2172
rect -11316 120 -7744 148
rect -7504 2172 -3932 2200
rect -7504 148 -4016 2172
rect -3952 148 -3932 2172
rect -7504 120 -3932 148
rect -3692 2172 -120 2200
rect -3692 148 -204 2172
rect -140 148 -120 2172
rect -3692 120 -120 148
rect 120 2172 3692 2200
rect 120 148 3608 2172
rect 3672 148 3692 2172
rect 120 120 3692 148
rect 3932 2172 7504 2200
rect 3932 148 7420 2172
rect 7484 148 7504 2172
rect 3932 120 7504 148
rect 7744 2172 11316 2200
rect 7744 148 11232 2172
rect 11296 148 11316 2172
rect 7744 120 11316 148
rect 11556 2172 15128 2200
rect 11556 148 15044 2172
rect 15108 148 15128 2172
rect 11556 120 15128 148
rect -15128 -148 -11556 -120
rect -15128 -2172 -11640 -148
rect -11576 -2172 -11556 -148
rect -15128 -2200 -11556 -2172
rect -11316 -148 -7744 -120
rect -11316 -2172 -7828 -148
rect -7764 -2172 -7744 -148
rect -11316 -2200 -7744 -2172
rect -7504 -148 -3932 -120
rect -7504 -2172 -4016 -148
rect -3952 -2172 -3932 -148
rect -7504 -2200 -3932 -2172
rect -3692 -148 -120 -120
rect -3692 -2172 -204 -148
rect -140 -2172 -120 -148
rect -3692 -2200 -120 -2172
rect 120 -148 3692 -120
rect 120 -2172 3608 -148
rect 3672 -2172 3692 -148
rect 120 -2200 3692 -2172
rect 3932 -148 7504 -120
rect 3932 -2172 7420 -148
rect 7484 -2172 7504 -148
rect 3932 -2200 7504 -2172
rect 7744 -148 11316 -120
rect 7744 -2172 11232 -148
rect 11296 -2172 11316 -148
rect 7744 -2200 11316 -2172
rect 11556 -148 15128 -120
rect 11556 -2172 15044 -148
rect 15108 -2172 15128 -148
rect 11556 -2200 15128 -2172
rect -15128 -2468 -11556 -2440
rect -15128 -4492 -11640 -2468
rect -11576 -4492 -11556 -2468
rect -15128 -4520 -11556 -4492
rect -11316 -2468 -7744 -2440
rect -11316 -4492 -7828 -2468
rect -7764 -4492 -7744 -2468
rect -11316 -4520 -7744 -4492
rect -7504 -2468 -3932 -2440
rect -7504 -4492 -4016 -2468
rect -3952 -4492 -3932 -2468
rect -7504 -4520 -3932 -4492
rect -3692 -2468 -120 -2440
rect -3692 -4492 -204 -2468
rect -140 -4492 -120 -2468
rect -3692 -4520 -120 -4492
rect 120 -2468 3692 -2440
rect 120 -4492 3608 -2468
rect 3672 -4492 3692 -2468
rect 120 -4520 3692 -4492
rect 3932 -2468 7504 -2440
rect 3932 -4492 7420 -2468
rect 7484 -4492 7504 -2468
rect 3932 -4520 7504 -4492
rect 7744 -2468 11316 -2440
rect 7744 -4492 11232 -2468
rect 11296 -4492 11316 -2468
rect 7744 -4520 11316 -4492
rect 11556 -2468 15128 -2440
rect 11556 -4492 15044 -2468
rect 15108 -4492 15128 -2468
rect 11556 -4520 15128 -4492
<< via3 >>
rect -11640 2468 -11576 4492
rect -7828 2468 -7764 4492
rect -4016 2468 -3952 4492
rect -204 2468 -140 4492
rect 3608 2468 3672 4492
rect 7420 2468 7484 4492
rect 11232 2468 11296 4492
rect 15044 2468 15108 4492
rect -11640 148 -11576 2172
rect -7828 148 -7764 2172
rect -4016 148 -3952 2172
rect -204 148 -140 2172
rect 3608 148 3672 2172
rect 7420 148 7484 2172
rect 11232 148 11296 2172
rect 15044 148 15108 2172
rect -11640 -2172 -11576 -148
rect -7828 -2172 -7764 -148
rect -4016 -2172 -3952 -148
rect -204 -2172 -140 -148
rect 3608 -2172 3672 -148
rect 7420 -2172 7484 -148
rect 11232 -2172 11296 -148
rect 15044 -2172 15108 -148
rect -11640 -4492 -11576 -2468
rect -7828 -4492 -7764 -2468
rect -4016 -4492 -3952 -2468
rect -204 -4492 -140 -2468
rect 3608 -4492 3672 -2468
rect 7420 -4492 7484 -2468
rect 11232 -4492 11296 -2468
rect 15044 -4492 15108 -2468
<< mimcap >>
rect -15088 4440 -11888 4480
rect -15088 2520 -15048 4440
rect -11928 2520 -11888 4440
rect -15088 2480 -11888 2520
rect -11276 4440 -8076 4480
rect -11276 2520 -11236 4440
rect -8116 2520 -8076 4440
rect -11276 2480 -8076 2520
rect -7464 4440 -4264 4480
rect -7464 2520 -7424 4440
rect -4304 2520 -4264 4440
rect -7464 2480 -4264 2520
rect -3652 4440 -452 4480
rect -3652 2520 -3612 4440
rect -492 2520 -452 4440
rect -3652 2480 -452 2520
rect 160 4440 3360 4480
rect 160 2520 200 4440
rect 3320 2520 3360 4440
rect 160 2480 3360 2520
rect 3972 4440 7172 4480
rect 3972 2520 4012 4440
rect 7132 2520 7172 4440
rect 3972 2480 7172 2520
rect 7784 4440 10984 4480
rect 7784 2520 7824 4440
rect 10944 2520 10984 4440
rect 7784 2480 10984 2520
rect 11596 4440 14796 4480
rect 11596 2520 11636 4440
rect 14756 2520 14796 4440
rect 11596 2480 14796 2520
rect -15088 2120 -11888 2160
rect -15088 200 -15048 2120
rect -11928 200 -11888 2120
rect -15088 160 -11888 200
rect -11276 2120 -8076 2160
rect -11276 200 -11236 2120
rect -8116 200 -8076 2120
rect -11276 160 -8076 200
rect -7464 2120 -4264 2160
rect -7464 200 -7424 2120
rect -4304 200 -4264 2120
rect -7464 160 -4264 200
rect -3652 2120 -452 2160
rect -3652 200 -3612 2120
rect -492 200 -452 2120
rect -3652 160 -452 200
rect 160 2120 3360 2160
rect 160 200 200 2120
rect 3320 200 3360 2120
rect 160 160 3360 200
rect 3972 2120 7172 2160
rect 3972 200 4012 2120
rect 7132 200 7172 2120
rect 3972 160 7172 200
rect 7784 2120 10984 2160
rect 7784 200 7824 2120
rect 10944 200 10984 2120
rect 7784 160 10984 200
rect 11596 2120 14796 2160
rect 11596 200 11636 2120
rect 14756 200 14796 2120
rect 11596 160 14796 200
rect -15088 -200 -11888 -160
rect -15088 -2120 -15048 -200
rect -11928 -2120 -11888 -200
rect -15088 -2160 -11888 -2120
rect -11276 -200 -8076 -160
rect -11276 -2120 -11236 -200
rect -8116 -2120 -8076 -200
rect -11276 -2160 -8076 -2120
rect -7464 -200 -4264 -160
rect -7464 -2120 -7424 -200
rect -4304 -2120 -4264 -200
rect -7464 -2160 -4264 -2120
rect -3652 -200 -452 -160
rect -3652 -2120 -3612 -200
rect -492 -2120 -452 -200
rect -3652 -2160 -452 -2120
rect 160 -200 3360 -160
rect 160 -2120 200 -200
rect 3320 -2120 3360 -200
rect 160 -2160 3360 -2120
rect 3972 -200 7172 -160
rect 3972 -2120 4012 -200
rect 7132 -2120 7172 -200
rect 3972 -2160 7172 -2120
rect 7784 -200 10984 -160
rect 7784 -2120 7824 -200
rect 10944 -2120 10984 -200
rect 7784 -2160 10984 -2120
rect 11596 -200 14796 -160
rect 11596 -2120 11636 -200
rect 14756 -2120 14796 -200
rect 11596 -2160 14796 -2120
rect -15088 -2520 -11888 -2480
rect -15088 -4440 -15048 -2520
rect -11928 -4440 -11888 -2520
rect -15088 -4480 -11888 -4440
rect -11276 -2520 -8076 -2480
rect -11276 -4440 -11236 -2520
rect -8116 -4440 -8076 -2520
rect -11276 -4480 -8076 -4440
rect -7464 -2520 -4264 -2480
rect -7464 -4440 -7424 -2520
rect -4304 -4440 -4264 -2520
rect -7464 -4480 -4264 -4440
rect -3652 -2520 -452 -2480
rect -3652 -4440 -3612 -2520
rect -492 -4440 -452 -2520
rect -3652 -4480 -452 -4440
rect 160 -2520 3360 -2480
rect 160 -4440 200 -2520
rect 3320 -4440 3360 -2520
rect 160 -4480 3360 -4440
rect 3972 -2520 7172 -2480
rect 3972 -4440 4012 -2520
rect 7132 -4440 7172 -2520
rect 3972 -4480 7172 -4440
rect 7784 -2520 10984 -2480
rect 7784 -4440 7824 -2520
rect 10944 -4440 10984 -2520
rect 7784 -4480 10984 -4440
rect 11596 -2520 14796 -2480
rect 11596 -4440 11636 -2520
rect 14756 -4440 14796 -2520
rect 11596 -4480 14796 -4440
<< mimcapcontact >>
rect -15048 2520 -11928 4440
rect -11236 2520 -8116 4440
rect -7424 2520 -4304 4440
rect -3612 2520 -492 4440
rect 200 2520 3320 4440
rect 4012 2520 7132 4440
rect 7824 2520 10944 4440
rect 11636 2520 14756 4440
rect -15048 200 -11928 2120
rect -11236 200 -8116 2120
rect -7424 200 -4304 2120
rect -3612 200 -492 2120
rect 200 200 3320 2120
rect 4012 200 7132 2120
rect 7824 200 10944 2120
rect 11636 200 14756 2120
rect -15048 -2120 -11928 -200
rect -11236 -2120 -8116 -200
rect -7424 -2120 -4304 -200
rect -3612 -2120 -492 -200
rect 200 -2120 3320 -200
rect 4012 -2120 7132 -200
rect 7824 -2120 10944 -200
rect 11636 -2120 14756 -200
rect -15048 -4440 -11928 -2520
rect -11236 -4440 -8116 -2520
rect -7424 -4440 -4304 -2520
rect -3612 -4440 -492 -2520
rect 200 -4440 3320 -2520
rect 4012 -4440 7132 -2520
rect 7824 -4440 10944 -2520
rect 11636 -4440 14756 -2520
<< metal4 >>
rect -11656 4492 -11560 4508
rect -15049 4440 -11927 4441
rect -15049 2520 -15048 4440
rect -11928 2520 -11927 4440
rect -15049 2519 -11927 2520
rect -11656 2468 -11640 4492
rect -11576 2468 -11560 4492
rect -7844 4492 -7748 4508
rect -11237 4440 -8115 4441
rect -11237 2520 -11236 4440
rect -8116 2520 -8115 4440
rect -11237 2519 -8115 2520
rect -11656 2452 -11560 2468
rect -7844 2468 -7828 4492
rect -7764 2468 -7748 4492
rect -4032 4492 -3936 4508
rect -7425 4440 -4303 4441
rect -7425 2520 -7424 4440
rect -4304 2520 -4303 4440
rect -7425 2519 -4303 2520
rect -7844 2452 -7748 2468
rect -4032 2468 -4016 4492
rect -3952 2468 -3936 4492
rect -220 4492 -124 4508
rect -3613 4440 -491 4441
rect -3613 2520 -3612 4440
rect -492 2520 -491 4440
rect -3613 2519 -491 2520
rect -4032 2452 -3936 2468
rect -220 2468 -204 4492
rect -140 2468 -124 4492
rect 3592 4492 3688 4508
rect 199 4440 3321 4441
rect 199 2520 200 4440
rect 3320 2520 3321 4440
rect 199 2519 3321 2520
rect -220 2452 -124 2468
rect 3592 2468 3608 4492
rect 3672 2468 3688 4492
rect 7404 4492 7500 4508
rect 4011 4440 7133 4441
rect 4011 2520 4012 4440
rect 7132 2520 7133 4440
rect 4011 2519 7133 2520
rect 3592 2452 3688 2468
rect 7404 2468 7420 4492
rect 7484 2468 7500 4492
rect 11216 4492 11312 4508
rect 7823 4440 10945 4441
rect 7823 2520 7824 4440
rect 10944 2520 10945 4440
rect 7823 2519 10945 2520
rect 7404 2452 7500 2468
rect 11216 2468 11232 4492
rect 11296 2468 11312 4492
rect 15028 4492 15124 4508
rect 11635 4440 14757 4441
rect 11635 2520 11636 4440
rect 14756 2520 14757 4440
rect 11635 2519 14757 2520
rect 11216 2452 11312 2468
rect 15028 2468 15044 4492
rect 15108 2468 15124 4492
rect 15028 2452 15124 2468
rect -11656 2172 -11560 2188
rect -15049 2120 -11927 2121
rect -15049 200 -15048 2120
rect -11928 200 -11927 2120
rect -15049 199 -11927 200
rect -11656 148 -11640 2172
rect -11576 148 -11560 2172
rect -7844 2172 -7748 2188
rect -11237 2120 -8115 2121
rect -11237 200 -11236 2120
rect -8116 200 -8115 2120
rect -11237 199 -8115 200
rect -11656 132 -11560 148
rect -7844 148 -7828 2172
rect -7764 148 -7748 2172
rect -4032 2172 -3936 2188
rect -7425 2120 -4303 2121
rect -7425 200 -7424 2120
rect -4304 200 -4303 2120
rect -7425 199 -4303 200
rect -7844 132 -7748 148
rect -4032 148 -4016 2172
rect -3952 148 -3936 2172
rect -220 2172 -124 2188
rect -3613 2120 -491 2121
rect -3613 200 -3612 2120
rect -492 200 -491 2120
rect -3613 199 -491 200
rect -4032 132 -3936 148
rect -220 148 -204 2172
rect -140 148 -124 2172
rect 3592 2172 3688 2188
rect 199 2120 3321 2121
rect 199 200 200 2120
rect 3320 200 3321 2120
rect 199 199 3321 200
rect -220 132 -124 148
rect 3592 148 3608 2172
rect 3672 148 3688 2172
rect 7404 2172 7500 2188
rect 4011 2120 7133 2121
rect 4011 200 4012 2120
rect 7132 200 7133 2120
rect 4011 199 7133 200
rect 3592 132 3688 148
rect 7404 148 7420 2172
rect 7484 148 7500 2172
rect 11216 2172 11312 2188
rect 7823 2120 10945 2121
rect 7823 200 7824 2120
rect 10944 200 10945 2120
rect 7823 199 10945 200
rect 7404 132 7500 148
rect 11216 148 11232 2172
rect 11296 148 11312 2172
rect 15028 2172 15124 2188
rect 11635 2120 14757 2121
rect 11635 200 11636 2120
rect 14756 200 14757 2120
rect 11635 199 14757 200
rect 11216 132 11312 148
rect 15028 148 15044 2172
rect 15108 148 15124 2172
rect 15028 132 15124 148
rect -11656 -148 -11560 -132
rect -15049 -200 -11927 -199
rect -15049 -2120 -15048 -200
rect -11928 -2120 -11927 -200
rect -15049 -2121 -11927 -2120
rect -11656 -2172 -11640 -148
rect -11576 -2172 -11560 -148
rect -7844 -148 -7748 -132
rect -11237 -200 -8115 -199
rect -11237 -2120 -11236 -200
rect -8116 -2120 -8115 -200
rect -11237 -2121 -8115 -2120
rect -11656 -2188 -11560 -2172
rect -7844 -2172 -7828 -148
rect -7764 -2172 -7748 -148
rect -4032 -148 -3936 -132
rect -7425 -200 -4303 -199
rect -7425 -2120 -7424 -200
rect -4304 -2120 -4303 -200
rect -7425 -2121 -4303 -2120
rect -7844 -2188 -7748 -2172
rect -4032 -2172 -4016 -148
rect -3952 -2172 -3936 -148
rect -220 -148 -124 -132
rect -3613 -200 -491 -199
rect -3613 -2120 -3612 -200
rect -492 -2120 -491 -200
rect -3613 -2121 -491 -2120
rect -4032 -2188 -3936 -2172
rect -220 -2172 -204 -148
rect -140 -2172 -124 -148
rect 3592 -148 3688 -132
rect 199 -200 3321 -199
rect 199 -2120 200 -200
rect 3320 -2120 3321 -200
rect 199 -2121 3321 -2120
rect -220 -2188 -124 -2172
rect 3592 -2172 3608 -148
rect 3672 -2172 3688 -148
rect 7404 -148 7500 -132
rect 4011 -200 7133 -199
rect 4011 -2120 4012 -200
rect 7132 -2120 7133 -200
rect 4011 -2121 7133 -2120
rect 3592 -2188 3688 -2172
rect 7404 -2172 7420 -148
rect 7484 -2172 7500 -148
rect 11216 -148 11312 -132
rect 7823 -200 10945 -199
rect 7823 -2120 7824 -200
rect 10944 -2120 10945 -200
rect 7823 -2121 10945 -2120
rect 7404 -2188 7500 -2172
rect 11216 -2172 11232 -148
rect 11296 -2172 11312 -148
rect 15028 -148 15124 -132
rect 11635 -200 14757 -199
rect 11635 -2120 11636 -200
rect 14756 -2120 14757 -200
rect 11635 -2121 14757 -2120
rect 11216 -2188 11312 -2172
rect 15028 -2172 15044 -148
rect 15108 -2172 15124 -148
rect 15028 -2188 15124 -2172
rect -11656 -2468 -11560 -2452
rect -15049 -2520 -11927 -2519
rect -15049 -4440 -15048 -2520
rect -11928 -4440 -11927 -2520
rect -15049 -4441 -11927 -4440
rect -11656 -4492 -11640 -2468
rect -11576 -4492 -11560 -2468
rect -7844 -2468 -7748 -2452
rect -11237 -2520 -8115 -2519
rect -11237 -4440 -11236 -2520
rect -8116 -4440 -8115 -2520
rect -11237 -4441 -8115 -4440
rect -11656 -4508 -11560 -4492
rect -7844 -4492 -7828 -2468
rect -7764 -4492 -7748 -2468
rect -4032 -2468 -3936 -2452
rect -7425 -2520 -4303 -2519
rect -7425 -4440 -7424 -2520
rect -4304 -4440 -4303 -2520
rect -7425 -4441 -4303 -4440
rect -7844 -4508 -7748 -4492
rect -4032 -4492 -4016 -2468
rect -3952 -4492 -3936 -2468
rect -220 -2468 -124 -2452
rect -3613 -2520 -491 -2519
rect -3613 -4440 -3612 -2520
rect -492 -4440 -491 -2520
rect -3613 -4441 -491 -4440
rect -4032 -4508 -3936 -4492
rect -220 -4492 -204 -2468
rect -140 -4492 -124 -2468
rect 3592 -2468 3688 -2452
rect 199 -2520 3321 -2519
rect 199 -4440 200 -2520
rect 3320 -4440 3321 -2520
rect 199 -4441 3321 -4440
rect -220 -4508 -124 -4492
rect 3592 -4492 3608 -2468
rect 3672 -4492 3688 -2468
rect 7404 -2468 7500 -2452
rect 4011 -2520 7133 -2519
rect 4011 -4440 4012 -2520
rect 7132 -4440 7133 -2520
rect 4011 -4441 7133 -4440
rect 3592 -4508 3688 -4492
rect 7404 -4492 7420 -2468
rect 7484 -4492 7500 -2468
rect 11216 -2468 11312 -2452
rect 7823 -2520 10945 -2519
rect 7823 -4440 7824 -2520
rect 10944 -4440 10945 -2520
rect 7823 -4441 10945 -4440
rect 7404 -4508 7500 -4492
rect 11216 -4492 11232 -2468
rect 11296 -4492 11312 -2468
rect 15028 -2468 15124 -2452
rect 11635 -2520 14757 -2519
rect 11635 -4440 11636 -2520
rect 14756 -4440 14757 -2520
rect 11635 -4441 14757 -4440
rect 11216 -4508 11312 -4492
rect 15028 -4492 15044 -2468
rect 15108 -4492 15124 -2468
rect 15028 -4508 15124 -4492
<< properties >>
string FIXED_BBOX 11556 2440 14836 4520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 16 l 10 val 329.88 carea 2.00 cperi 0.19 nx 8 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>

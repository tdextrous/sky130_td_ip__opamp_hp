magic
tech sky130A
magscale 1 2
timestamp 1713233716
<< nwell >>
rect -2293 -497 2293 497
<< mvpmos >>
rect -2035 -200 -1835 200
rect -1777 -200 -1577 200
rect -1519 -200 -1319 200
rect -1261 -200 -1061 200
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
rect 1061 -200 1261 200
rect 1319 -200 1519 200
rect 1577 -200 1777 200
rect 1835 -200 2035 200
<< mvpdiff >>
rect -2093 188 -2035 200
rect -2093 -188 -2081 188
rect -2047 -188 -2035 188
rect -2093 -200 -2035 -188
rect -1835 188 -1777 200
rect -1835 -188 -1823 188
rect -1789 -188 -1777 188
rect -1835 -200 -1777 -188
rect -1577 188 -1519 200
rect -1577 -188 -1565 188
rect -1531 -188 -1519 188
rect -1577 -200 -1519 -188
rect -1319 188 -1261 200
rect -1319 -188 -1307 188
rect -1273 -188 -1261 188
rect -1319 -200 -1261 -188
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
rect 1261 188 1319 200
rect 1261 -188 1273 188
rect 1307 -188 1319 188
rect 1261 -200 1319 -188
rect 1519 188 1577 200
rect 1519 -188 1531 188
rect 1565 -188 1577 188
rect 1519 -200 1577 -188
rect 1777 188 1835 200
rect 1777 -188 1789 188
rect 1823 -188 1835 188
rect 1777 -200 1835 -188
rect 2035 188 2093 200
rect 2035 -188 2047 188
rect 2081 -188 2093 188
rect 2035 -200 2093 -188
<< mvpdiffc >>
rect -2081 -188 -2047 188
rect -1823 -188 -1789 188
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect 1789 -188 1823 188
rect 2047 -188 2081 188
<< mvnsubdiff >>
rect -2227 419 2227 431
rect -2227 385 -2119 419
rect 2119 385 2227 419
rect -2227 373 2227 385
rect -2227 323 -2169 373
rect -2227 -323 -2215 323
rect -2181 -323 -2169 323
rect 2169 323 2227 373
rect -2227 -373 -2169 -323
rect 2169 -323 2181 323
rect 2215 -323 2227 323
rect 2169 -373 2227 -323
rect -2227 -385 2227 -373
rect -2227 -419 -2119 -385
rect 2119 -419 2227 -385
rect -2227 -431 2227 -419
<< mvnsubdiffcont >>
rect -2119 385 2119 419
rect -2215 -323 -2181 323
rect 2181 -323 2215 323
rect -2119 -419 2119 -385
<< poly >>
rect -2035 281 -1835 297
rect -2035 247 -2019 281
rect -1851 247 -1835 281
rect -2035 200 -1835 247
rect -1777 281 -1577 297
rect -1777 247 -1761 281
rect -1593 247 -1577 281
rect -1777 200 -1577 247
rect -1519 281 -1319 297
rect -1519 247 -1503 281
rect -1335 247 -1319 281
rect -1519 200 -1319 247
rect -1261 281 -1061 297
rect -1261 247 -1245 281
rect -1077 247 -1061 281
rect -1261 200 -1061 247
rect -1003 281 -803 297
rect -1003 247 -987 281
rect -819 247 -803 281
rect -1003 200 -803 247
rect -745 281 -545 297
rect -745 247 -729 281
rect -561 247 -545 281
rect -745 200 -545 247
rect -487 281 -287 297
rect -487 247 -471 281
rect -303 247 -287 281
rect -487 200 -287 247
rect -229 281 -29 297
rect -229 247 -213 281
rect -45 247 -29 281
rect -229 200 -29 247
rect 29 281 229 297
rect 29 247 45 281
rect 213 247 229 281
rect 29 200 229 247
rect 287 281 487 297
rect 287 247 303 281
rect 471 247 487 281
rect 287 200 487 247
rect 545 281 745 297
rect 545 247 561 281
rect 729 247 745 281
rect 545 200 745 247
rect 803 281 1003 297
rect 803 247 819 281
rect 987 247 1003 281
rect 803 200 1003 247
rect 1061 281 1261 297
rect 1061 247 1077 281
rect 1245 247 1261 281
rect 1061 200 1261 247
rect 1319 281 1519 297
rect 1319 247 1335 281
rect 1503 247 1519 281
rect 1319 200 1519 247
rect 1577 281 1777 297
rect 1577 247 1593 281
rect 1761 247 1777 281
rect 1577 200 1777 247
rect 1835 281 2035 297
rect 1835 247 1851 281
rect 2019 247 2035 281
rect 1835 200 2035 247
rect -2035 -247 -1835 -200
rect -2035 -281 -2019 -247
rect -1851 -281 -1835 -247
rect -2035 -297 -1835 -281
rect -1777 -247 -1577 -200
rect -1777 -281 -1761 -247
rect -1593 -281 -1577 -247
rect -1777 -297 -1577 -281
rect -1519 -247 -1319 -200
rect -1519 -281 -1503 -247
rect -1335 -281 -1319 -247
rect -1519 -297 -1319 -281
rect -1261 -247 -1061 -200
rect -1261 -281 -1245 -247
rect -1077 -281 -1061 -247
rect -1261 -297 -1061 -281
rect -1003 -247 -803 -200
rect -1003 -281 -987 -247
rect -819 -281 -803 -247
rect -1003 -297 -803 -281
rect -745 -247 -545 -200
rect -745 -281 -729 -247
rect -561 -281 -545 -247
rect -745 -297 -545 -281
rect -487 -247 -287 -200
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -487 -297 -287 -281
rect -229 -247 -29 -200
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect -229 -297 -29 -281
rect 29 -247 229 -200
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 29 -297 229 -281
rect 287 -247 487 -200
rect 287 -281 303 -247
rect 471 -281 487 -247
rect 287 -297 487 -281
rect 545 -247 745 -200
rect 545 -281 561 -247
rect 729 -281 745 -247
rect 545 -297 745 -281
rect 803 -247 1003 -200
rect 803 -281 819 -247
rect 987 -281 1003 -247
rect 803 -297 1003 -281
rect 1061 -247 1261 -200
rect 1061 -281 1077 -247
rect 1245 -281 1261 -247
rect 1061 -297 1261 -281
rect 1319 -247 1519 -200
rect 1319 -281 1335 -247
rect 1503 -281 1519 -247
rect 1319 -297 1519 -281
rect 1577 -247 1777 -200
rect 1577 -281 1593 -247
rect 1761 -281 1777 -247
rect 1577 -297 1777 -281
rect 1835 -247 2035 -200
rect 1835 -281 1851 -247
rect 2019 -281 2035 -247
rect 1835 -297 2035 -281
<< polycont >>
rect -2019 247 -1851 281
rect -1761 247 -1593 281
rect -1503 247 -1335 281
rect -1245 247 -1077 281
rect -987 247 -819 281
rect -729 247 -561 281
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect 561 247 729 281
rect 819 247 987 281
rect 1077 247 1245 281
rect 1335 247 1503 281
rect 1593 247 1761 281
rect 1851 247 2019 281
rect -2019 -281 -1851 -247
rect -1761 -281 -1593 -247
rect -1503 -281 -1335 -247
rect -1245 -281 -1077 -247
rect -987 -281 -819 -247
rect -729 -281 -561 -247
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
rect 561 -281 729 -247
rect 819 -281 987 -247
rect 1077 -281 1245 -247
rect 1335 -281 1503 -247
rect 1593 -281 1761 -247
rect 1851 -281 2019 -247
<< locali >>
rect -2215 385 -2119 419
rect 2119 385 2215 419
rect -2215 323 -2181 385
rect 2181 323 2215 385
rect -2035 247 -2019 281
rect -1851 247 -1835 281
rect -1777 247 -1761 281
rect -1593 247 -1577 281
rect -1519 247 -1503 281
rect -1335 247 -1319 281
rect -1261 247 -1245 281
rect -1077 247 -1061 281
rect -1003 247 -987 281
rect -819 247 -803 281
rect -745 247 -729 281
rect -561 247 -545 281
rect -487 247 -471 281
rect -303 247 -287 281
rect -229 247 -213 281
rect -45 247 -29 281
rect 29 247 45 281
rect 213 247 229 281
rect 287 247 303 281
rect 471 247 487 281
rect 545 247 561 281
rect 729 247 745 281
rect 803 247 819 281
rect 987 247 1003 281
rect 1061 247 1077 281
rect 1245 247 1261 281
rect 1319 247 1335 281
rect 1503 247 1519 281
rect 1577 247 1593 281
rect 1761 247 1777 281
rect 1835 247 1851 281
rect 2019 247 2035 281
rect -2081 188 -2047 204
rect -2081 -204 -2047 -188
rect -1823 188 -1789 204
rect -1823 -204 -1789 -188
rect -1565 188 -1531 204
rect -1565 -204 -1531 -188
rect -1307 188 -1273 204
rect -1307 -204 -1273 -188
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect 1273 188 1307 204
rect 1273 -204 1307 -188
rect 1531 188 1565 204
rect 1531 -204 1565 -188
rect 1789 188 1823 204
rect 1789 -204 1823 -188
rect 2047 188 2081 204
rect 2047 -204 2081 -188
rect -2035 -281 -2019 -247
rect -1851 -281 -1835 -247
rect -1777 -281 -1761 -247
rect -1593 -281 -1577 -247
rect -1519 -281 -1503 -247
rect -1335 -281 -1319 -247
rect -1261 -281 -1245 -247
rect -1077 -281 -1061 -247
rect -1003 -281 -987 -247
rect -819 -281 -803 -247
rect -745 -281 -729 -247
rect -561 -281 -545 -247
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 287 -281 303 -247
rect 471 -281 487 -247
rect 545 -281 561 -247
rect 729 -281 745 -247
rect 803 -281 819 -247
rect 987 -281 1003 -247
rect 1061 -281 1077 -247
rect 1245 -281 1261 -247
rect 1319 -281 1335 -247
rect 1503 -281 1519 -247
rect 1577 -281 1593 -247
rect 1761 -281 1777 -247
rect 1835 -281 1851 -247
rect 2019 -281 2035 -247
rect -2215 -385 -2181 -323
rect 2181 -385 2215 -323
rect -2215 -419 -2119 -385
rect 2119 -419 2215 -385
<< viali >>
rect -2019 247 -1851 281
rect -1761 247 -1593 281
rect -1503 247 -1335 281
rect -1245 247 -1077 281
rect -987 247 -819 281
rect -729 247 -561 281
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect 561 247 729 281
rect 819 247 987 281
rect 1077 247 1245 281
rect 1335 247 1503 281
rect 1593 247 1761 281
rect 1851 247 2019 281
rect -2081 -188 -2047 188
rect -1823 -188 -1789 188
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect 1789 -188 1823 188
rect 2047 -188 2081 188
rect -2019 -281 -1851 -247
rect -1761 -281 -1593 -247
rect -1503 -281 -1335 -247
rect -1245 -281 -1077 -247
rect -987 -281 -819 -247
rect -729 -281 -561 -247
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
rect 561 -281 729 -247
rect 819 -281 987 -247
rect 1077 -281 1245 -247
rect 1335 -281 1503 -247
rect 1593 -281 1761 -247
rect 1851 -281 2019 -247
<< metal1 >>
rect -2031 281 -1839 287
rect -2031 247 -2019 281
rect -1851 247 -1839 281
rect -2031 241 -1839 247
rect -1773 281 -1581 287
rect -1773 247 -1761 281
rect -1593 247 -1581 281
rect -1773 241 -1581 247
rect -1515 281 -1323 287
rect -1515 247 -1503 281
rect -1335 247 -1323 281
rect -1515 241 -1323 247
rect -1257 281 -1065 287
rect -1257 247 -1245 281
rect -1077 247 -1065 281
rect -1257 241 -1065 247
rect -999 281 -807 287
rect -999 247 -987 281
rect -819 247 -807 281
rect -999 241 -807 247
rect -741 281 -549 287
rect -741 247 -729 281
rect -561 247 -549 281
rect -741 241 -549 247
rect -483 281 -291 287
rect -483 247 -471 281
rect -303 247 -291 281
rect -483 241 -291 247
rect -225 281 -33 287
rect -225 247 -213 281
rect -45 247 -33 281
rect -225 241 -33 247
rect 33 281 225 287
rect 33 247 45 281
rect 213 247 225 281
rect 33 241 225 247
rect 291 281 483 287
rect 291 247 303 281
rect 471 247 483 281
rect 291 241 483 247
rect 549 281 741 287
rect 549 247 561 281
rect 729 247 741 281
rect 549 241 741 247
rect 807 281 999 287
rect 807 247 819 281
rect 987 247 999 281
rect 807 241 999 247
rect 1065 281 1257 287
rect 1065 247 1077 281
rect 1245 247 1257 281
rect 1065 241 1257 247
rect 1323 281 1515 287
rect 1323 247 1335 281
rect 1503 247 1515 281
rect 1323 241 1515 247
rect 1581 281 1773 287
rect 1581 247 1593 281
rect 1761 247 1773 281
rect 1581 241 1773 247
rect 1839 281 2031 287
rect 1839 247 1851 281
rect 2019 247 2031 281
rect 1839 241 2031 247
rect -2087 188 -2041 200
rect -2087 -188 -2081 188
rect -2047 -188 -2041 188
rect -2087 -200 -2041 -188
rect -1829 188 -1783 200
rect -1829 -188 -1823 188
rect -1789 -188 -1783 188
rect -1829 -200 -1783 -188
rect -1571 188 -1525 200
rect -1571 -188 -1565 188
rect -1531 -188 -1525 188
rect -1571 -200 -1525 -188
rect -1313 188 -1267 200
rect -1313 -188 -1307 188
rect -1273 -188 -1267 188
rect -1313 -200 -1267 -188
rect -1055 188 -1009 200
rect -1055 -188 -1049 188
rect -1015 -188 -1009 188
rect -1055 -200 -1009 -188
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect 1009 188 1055 200
rect 1009 -188 1015 188
rect 1049 -188 1055 188
rect 1009 -200 1055 -188
rect 1267 188 1313 200
rect 1267 -188 1273 188
rect 1307 -188 1313 188
rect 1267 -200 1313 -188
rect 1525 188 1571 200
rect 1525 -188 1531 188
rect 1565 -188 1571 188
rect 1525 -200 1571 -188
rect 1783 188 1829 200
rect 1783 -188 1789 188
rect 1823 -188 1829 188
rect 1783 -200 1829 -188
rect 2041 188 2087 200
rect 2041 -188 2047 188
rect 2081 -188 2087 188
rect 2041 -200 2087 -188
rect -2031 -247 -1839 -241
rect -2031 -281 -2019 -247
rect -1851 -281 -1839 -247
rect -2031 -287 -1839 -281
rect -1773 -247 -1581 -241
rect -1773 -281 -1761 -247
rect -1593 -281 -1581 -247
rect -1773 -287 -1581 -281
rect -1515 -247 -1323 -241
rect -1515 -281 -1503 -247
rect -1335 -281 -1323 -247
rect -1515 -287 -1323 -281
rect -1257 -247 -1065 -241
rect -1257 -281 -1245 -247
rect -1077 -281 -1065 -247
rect -1257 -287 -1065 -281
rect -999 -247 -807 -241
rect -999 -281 -987 -247
rect -819 -281 -807 -247
rect -999 -287 -807 -281
rect -741 -247 -549 -241
rect -741 -281 -729 -247
rect -561 -281 -549 -247
rect -741 -287 -549 -281
rect -483 -247 -291 -241
rect -483 -281 -471 -247
rect -303 -281 -291 -247
rect -483 -287 -291 -281
rect -225 -247 -33 -241
rect -225 -281 -213 -247
rect -45 -281 -33 -247
rect -225 -287 -33 -281
rect 33 -247 225 -241
rect 33 -281 45 -247
rect 213 -281 225 -247
rect 33 -287 225 -281
rect 291 -247 483 -241
rect 291 -281 303 -247
rect 471 -281 483 -247
rect 291 -287 483 -281
rect 549 -247 741 -241
rect 549 -281 561 -247
rect 729 -281 741 -247
rect 549 -287 741 -281
rect 807 -247 999 -241
rect 807 -281 819 -247
rect 987 -281 999 -247
rect 807 -287 999 -281
rect 1065 -247 1257 -241
rect 1065 -281 1077 -247
rect 1245 -281 1257 -247
rect 1065 -287 1257 -281
rect 1323 -247 1515 -241
rect 1323 -281 1335 -247
rect 1503 -281 1515 -247
rect 1323 -287 1515 -281
rect 1581 -247 1773 -241
rect 1581 -281 1593 -247
rect 1761 -281 1773 -247
rect 1581 -287 1773 -281
rect 1839 -247 2031 -241
rect 1839 -281 1851 -247
rect 2019 -281 2031 -247
rect 1839 -287 2031 -281
<< properties >>
string FIXED_BBOX -2198 -402 2198 402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

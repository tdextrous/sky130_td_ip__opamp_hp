magic
tech sky130A
magscale 1 2
timestamp 1713674343
<< pwell >>
rect -586 -722 586 722
<< psubdiff >>
rect -550 652 -454 686
rect 454 652 550 686
rect -550 590 -516 652
rect 516 590 550 652
rect -550 -652 -516 -590
rect 516 -652 550 -590
rect -550 -686 -454 -652
rect 454 -686 550 -652
<< psubdiffcont >>
rect -454 652 454 686
rect -550 -590 -516 590
rect 516 -590 550 590
rect -454 -686 454 -652
<< xpolycontact >>
rect -420 124 -282 556
rect -420 -556 -282 -124
rect -186 124 -48 556
rect -186 -556 -48 -124
rect 48 124 186 556
rect 48 -556 186 -124
rect 282 124 420 556
rect 282 -556 420 -124
<< ppolyres >>
rect -420 -124 -282 124
rect -186 -124 -48 124
rect 48 -124 186 124
rect 282 -124 420 124
<< locali >>
rect -550 652 -454 686
rect 454 652 550 686
rect -550 590 -516 652
rect 516 590 550 652
rect -550 -652 -516 -590
rect 516 -652 550 -590
rect -550 -686 -454 -652
rect 454 -686 550 -652
<< viali >>
rect -404 141 -298 538
rect -170 141 -64 538
rect 64 141 170 538
rect 298 141 404 538
rect -404 -538 -298 -141
rect -170 -538 -64 -141
rect 64 -538 170 -141
rect 298 -538 404 -141
<< metal1 >>
rect -410 538 -292 550
rect -410 141 -404 538
rect -298 141 -292 538
rect -410 129 -292 141
rect -176 538 -58 550
rect -176 141 -170 538
rect -64 141 -58 538
rect -176 129 -58 141
rect 58 538 176 550
rect 58 141 64 538
rect 170 141 176 538
rect 58 129 176 141
rect 292 538 410 550
rect 292 141 298 538
rect 404 141 410 538
rect 292 129 410 141
rect -410 -141 -292 -129
rect -410 -538 -404 -141
rect -298 -538 -292 -141
rect -410 -550 -292 -538
rect -176 -141 -58 -129
rect -176 -538 -170 -141
rect -64 -538 -58 -141
rect -176 -550 -58 -538
rect 58 -141 176 -129
rect 58 -538 64 -141
rect 170 -538 176 -141
rect 58 -550 176 -538
rect 292 -141 410 -129
rect 292 -538 298 -141
rect 404 -538 410 -141
rect 292 -550 410 -538
<< properties >>
string FIXED_BBOX -533 -669 533 669
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 1.4 m 1 nx 4 wmin 0.690 lmin 0.50 rho 319.8 val 1.213k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713306471
<< pwell >>
rect -3553 -558 3553 558
<< mvnmos >>
rect -3325 -300 -3125 300
rect -3067 -300 -2867 300
rect -2809 -300 -2609 300
rect -2551 -300 -2351 300
rect -2293 -300 -2093 300
rect -2035 -300 -1835 300
rect -1777 -300 -1577 300
rect -1519 -300 -1319 300
rect -1261 -300 -1061 300
rect -1003 -300 -803 300
rect -745 -300 -545 300
rect -487 -300 -287 300
rect -229 -300 -29 300
rect 29 -300 229 300
rect 287 -300 487 300
rect 545 -300 745 300
rect 803 -300 1003 300
rect 1061 -300 1261 300
rect 1319 -300 1519 300
rect 1577 -300 1777 300
rect 1835 -300 2035 300
rect 2093 -300 2293 300
rect 2351 -300 2551 300
rect 2609 -300 2809 300
rect 2867 -300 3067 300
rect 3125 -300 3325 300
<< mvndiff >>
rect -3383 288 -3325 300
rect -3383 -288 -3371 288
rect -3337 -288 -3325 288
rect -3383 -300 -3325 -288
rect -3125 288 -3067 300
rect -3125 -288 -3113 288
rect -3079 -288 -3067 288
rect -3125 -300 -3067 -288
rect -2867 288 -2809 300
rect -2867 -288 -2855 288
rect -2821 -288 -2809 288
rect -2867 -300 -2809 -288
rect -2609 288 -2551 300
rect -2609 -288 -2597 288
rect -2563 -288 -2551 288
rect -2609 -300 -2551 -288
rect -2351 288 -2293 300
rect -2351 -288 -2339 288
rect -2305 -288 -2293 288
rect -2351 -300 -2293 -288
rect -2093 288 -2035 300
rect -2093 -288 -2081 288
rect -2047 -288 -2035 288
rect -2093 -300 -2035 -288
rect -1835 288 -1777 300
rect -1835 -288 -1823 288
rect -1789 -288 -1777 288
rect -1835 -300 -1777 -288
rect -1577 288 -1519 300
rect -1577 -288 -1565 288
rect -1531 -288 -1519 288
rect -1577 -300 -1519 -288
rect -1319 288 -1261 300
rect -1319 -288 -1307 288
rect -1273 -288 -1261 288
rect -1319 -300 -1261 -288
rect -1061 288 -1003 300
rect -1061 -288 -1049 288
rect -1015 -288 -1003 288
rect -1061 -300 -1003 -288
rect -803 288 -745 300
rect -803 -288 -791 288
rect -757 -288 -745 288
rect -803 -300 -745 -288
rect -545 288 -487 300
rect -545 -288 -533 288
rect -499 -288 -487 288
rect -545 -300 -487 -288
rect -287 288 -229 300
rect -287 -288 -275 288
rect -241 -288 -229 288
rect -287 -300 -229 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 229 288 287 300
rect 229 -288 241 288
rect 275 -288 287 288
rect 229 -300 287 -288
rect 487 288 545 300
rect 487 -288 499 288
rect 533 -288 545 288
rect 487 -300 545 -288
rect 745 288 803 300
rect 745 -288 757 288
rect 791 -288 803 288
rect 745 -300 803 -288
rect 1003 288 1061 300
rect 1003 -288 1015 288
rect 1049 -288 1061 288
rect 1003 -300 1061 -288
rect 1261 288 1319 300
rect 1261 -288 1273 288
rect 1307 -288 1319 288
rect 1261 -300 1319 -288
rect 1519 288 1577 300
rect 1519 -288 1531 288
rect 1565 -288 1577 288
rect 1519 -300 1577 -288
rect 1777 288 1835 300
rect 1777 -288 1789 288
rect 1823 -288 1835 288
rect 1777 -300 1835 -288
rect 2035 288 2093 300
rect 2035 -288 2047 288
rect 2081 -288 2093 288
rect 2035 -300 2093 -288
rect 2293 288 2351 300
rect 2293 -288 2305 288
rect 2339 -288 2351 288
rect 2293 -300 2351 -288
rect 2551 288 2609 300
rect 2551 -288 2563 288
rect 2597 -288 2609 288
rect 2551 -300 2609 -288
rect 2809 288 2867 300
rect 2809 -288 2821 288
rect 2855 -288 2867 288
rect 2809 -300 2867 -288
rect 3067 288 3125 300
rect 3067 -288 3079 288
rect 3113 -288 3125 288
rect 3067 -300 3125 -288
rect 3325 288 3383 300
rect 3325 -288 3337 288
rect 3371 -288 3383 288
rect 3325 -300 3383 -288
<< mvndiffc >>
rect -3371 -288 -3337 288
rect -3113 -288 -3079 288
rect -2855 -288 -2821 288
rect -2597 -288 -2563 288
rect -2339 -288 -2305 288
rect -2081 -288 -2047 288
rect -1823 -288 -1789 288
rect -1565 -288 -1531 288
rect -1307 -288 -1273 288
rect -1049 -288 -1015 288
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect 1015 -288 1049 288
rect 1273 -288 1307 288
rect 1531 -288 1565 288
rect 1789 -288 1823 288
rect 2047 -288 2081 288
rect 2305 -288 2339 288
rect 2563 -288 2597 288
rect 2821 -288 2855 288
rect 3079 -288 3113 288
rect 3337 -288 3371 288
<< mvpsubdiff >>
rect -3517 510 3517 522
rect -3517 476 -3409 510
rect 3409 476 3517 510
rect -3517 464 3517 476
rect -3517 414 -3459 464
rect -3517 -414 -3505 414
rect -3471 -414 -3459 414
rect 3459 414 3517 464
rect -3517 -464 -3459 -414
rect 3459 -414 3471 414
rect 3505 -414 3517 414
rect 3459 -464 3517 -414
rect -3517 -476 3517 -464
rect -3517 -510 -3409 -476
rect 3409 -510 3517 -476
rect -3517 -522 3517 -510
<< mvpsubdiffcont >>
rect -3409 476 3409 510
rect -3505 -414 -3471 414
rect 3471 -414 3505 414
rect -3409 -510 3409 -476
<< poly >>
rect -3291 372 -3159 388
rect -3291 355 -3275 372
rect -3325 338 -3275 355
rect -3175 355 -3159 372
rect -3033 372 -2901 388
rect -3033 355 -3017 372
rect -3175 338 -3125 355
rect -3325 300 -3125 338
rect -3067 338 -3017 355
rect -2917 355 -2901 372
rect -2775 372 -2643 388
rect -2775 355 -2759 372
rect -2917 338 -2867 355
rect -3067 300 -2867 338
rect -2809 338 -2759 355
rect -2659 355 -2643 372
rect -2517 372 -2385 388
rect -2517 355 -2501 372
rect -2659 338 -2609 355
rect -2809 300 -2609 338
rect -2551 338 -2501 355
rect -2401 355 -2385 372
rect -2259 372 -2127 388
rect -2259 355 -2243 372
rect -2401 338 -2351 355
rect -2551 300 -2351 338
rect -2293 338 -2243 355
rect -2143 355 -2127 372
rect -2001 372 -1869 388
rect -2001 355 -1985 372
rect -2143 338 -2093 355
rect -2293 300 -2093 338
rect -2035 338 -1985 355
rect -1885 355 -1869 372
rect -1743 372 -1611 388
rect -1743 355 -1727 372
rect -1885 338 -1835 355
rect -2035 300 -1835 338
rect -1777 338 -1727 355
rect -1627 355 -1611 372
rect -1485 372 -1353 388
rect -1485 355 -1469 372
rect -1627 338 -1577 355
rect -1777 300 -1577 338
rect -1519 338 -1469 355
rect -1369 355 -1353 372
rect -1227 372 -1095 388
rect -1227 355 -1211 372
rect -1369 338 -1319 355
rect -1519 300 -1319 338
rect -1261 338 -1211 355
rect -1111 355 -1095 372
rect -969 372 -837 388
rect -969 355 -953 372
rect -1111 338 -1061 355
rect -1261 300 -1061 338
rect -1003 338 -953 355
rect -853 355 -837 372
rect -711 372 -579 388
rect -711 355 -695 372
rect -853 338 -803 355
rect -1003 300 -803 338
rect -745 338 -695 355
rect -595 355 -579 372
rect -453 372 -321 388
rect -453 355 -437 372
rect -595 338 -545 355
rect -745 300 -545 338
rect -487 338 -437 355
rect -337 355 -321 372
rect -195 372 -63 388
rect -195 355 -179 372
rect -337 338 -287 355
rect -487 300 -287 338
rect -229 338 -179 355
rect -79 355 -63 372
rect 63 372 195 388
rect 63 355 79 372
rect -79 338 -29 355
rect -229 300 -29 338
rect 29 338 79 355
rect 179 355 195 372
rect 321 372 453 388
rect 321 355 337 372
rect 179 338 229 355
rect 29 300 229 338
rect 287 338 337 355
rect 437 355 453 372
rect 579 372 711 388
rect 579 355 595 372
rect 437 338 487 355
rect 287 300 487 338
rect 545 338 595 355
rect 695 355 711 372
rect 837 372 969 388
rect 837 355 853 372
rect 695 338 745 355
rect 545 300 745 338
rect 803 338 853 355
rect 953 355 969 372
rect 1095 372 1227 388
rect 1095 355 1111 372
rect 953 338 1003 355
rect 803 300 1003 338
rect 1061 338 1111 355
rect 1211 355 1227 372
rect 1353 372 1485 388
rect 1353 355 1369 372
rect 1211 338 1261 355
rect 1061 300 1261 338
rect 1319 338 1369 355
rect 1469 355 1485 372
rect 1611 372 1743 388
rect 1611 355 1627 372
rect 1469 338 1519 355
rect 1319 300 1519 338
rect 1577 338 1627 355
rect 1727 355 1743 372
rect 1869 372 2001 388
rect 1869 355 1885 372
rect 1727 338 1777 355
rect 1577 300 1777 338
rect 1835 338 1885 355
rect 1985 355 2001 372
rect 2127 372 2259 388
rect 2127 355 2143 372
rect 1985 338 2035 355
rect 1835 300 2035 338
rect 2093 338 2143 355
rect 2243 355 2259 372
rect 2385 372 2517 388
rect 2385 355 2401 372
rect 2243 338 2293 355
rect 2093 300 2293 338
rect 2351 338 2401 355
rect 2501 355 2517 372
rect 2643 372 2775 388
rect 2643 355 2659 372
rect 2501 338 2551 355
rect 2351 300 2551 338
rect 2609 338 2659 355
rect 2759 355 2775 372
rect 2901 372 3033 388
rect 2901 355 2917 372
rect 2759 338 2809 355
rect 2609 300 2809 338
rect 2867 338 2917 355
rect 3017 355 3033 372
rect 3159 372 3291 388
rect 3159 355 3175 372
rect 3017 338 3067 355
rect 2867 300 3067 338
rect 3125 338 3175 355
rect 3275 355 3291 372
rect 3275 338 3325 355
rect 3125 300 3325 338
rect -3325 -338 -3125 -300
rect -3325 -355 -3275 -338
rect -3291 -372 -3275 -355
rect -3175 -355 -3125 -338
rect -3067 -338 -2867 -300
rect -3067 -355 -3017 -338
rect -3175 -372 -3159 -355
rect -3291 -388 -3159 -372
rect -3033 -372 -3017 -355
rect -2917 -355 -2867 -338
rect -2809 -338 -2609 -300
rect -2809 -355 -2759 -338
rect -2917 -372 -2901 -355
rect -3033 -388 -2901 -372
rect -2775 -372 -2759 -355
rect -2659 -355 -2609 -338
rect -2551 -338 -2351 -300
rect -2551 -355 -2501 -338
rect -2659 -372 -2643 -355
rect -2775 -388 -2643 -372
rect -2517 -372 -2501 -355
rect -2401 -355 -2351 -338
rect -2293 -338 -2093 -300
rect -2293 -355 -2243 -338
rect -2401 -372 -2385 -355
rect -2517 -388 -2385 -372
rect -2259 -372 -2243 -355
rect -2143 -355 -2093 -338
rect -2035 -338 -1835 -300
rect -2035 -355 -1985 -338
rect -2143 -372 -2127 -355
rect -2259 -388 -2127 -372
rect -2001 -372 -1985 -355
rect -1885 -355 -1835 -338
rect -1777 -338 -1577 -300
rect -1777 -355 -1727 -338
rect -1885 -372 -1869 -355
rect -2001 -388 -1869 -372
rect -1743 -372 -1727 -355
rect -1627 -355 -1577 -338
rect -1519 -338 -1319 -300
rect -1519 -355 -1469 -338
rect -1627 -372 -1611 -355
rect -1743 -388 -1611 -372
rect -1485 -372 -1469 -355
rect -1369 -355 -1319 -338
rect -1261 -338 -1061 -300
rect -1261 -355 -1211 -338
rect -1369 -372 -1353 -355
rect -1485 -388 -1353 -372
rect -1227 -372 -1211 -355
rect -1111 -355 -1061 -338
rect -1003 -338 -803 -300
rect -1003 -355 -953 -338
rect -1111 -372 -1095 -355
rect -1227 -388 -1095 -372
rect -969 -372 -953 -355
rect -853 -355 -803 -338
rect -745 -338 -545 -300
rect -745 -355 -695 -338
rect -853 -372 -837 -355
rect -969 -388 -837 -372
rect -711 -372 -695 -355
rect -595 -355 -545 -338
rect -487 -338 -287 -300
rect -487 -355 -437 -338
rect -595 -372 -579 -355
rect -711 -388 -579 -372
rect -453 -372 -437 -355
rect -337 -355 -287 -338
rect -229 -338 -29 -300
rect -229 -355 -179 -338
rect -337 -372 -321 -355
rect -453 -388 -321 -372
rect -195 -372 -179 -355
rect -79 -355 -29 -338
rect 29 -338 229 -300
rect 29 -355 79 -338
rect -79 -372 -63 -355
rect -195 -388 -63 -372
rect 63 -372 79 -355
rect 179 -355 229 -338
rect 287 -338 487 -300
rect 287 -355 337 -338
rect 179 -372 195 -355
rect 63 -388 195 -372
rect 321 -372 337 -355
rect 437 -355 487 -338
rect 545 -338 745 -300
rect 545 -355 595 -338
rect 437 -372 453 -355
rect 321 -388 453 -372
rect 579 -372 595 -355
rect 695 -355 745 -338
rect 803 -338 1003 -300
rect 803 -355 853 -338
rect 695 -372 711 -355
rect 579 -388 711 -372
rect 837 -372 853 -355
rect 953 -355 1003 -338
rect 1061 -338 1261 -300
rect 1061 -355 1111 -338
rect 953 -372 969 -355
rect 837 -388 969 -372
rect 1095 -372 1111 -355
rect 1211 -355 1261 -338
rect 1319 -338 1519 -300
rect 1319 -355 1369 -338
rect 1211 -372 1227 -355
rect 1095 -388 1227 -372
rect 1353 -372 1369 -355
rect 1469 -355 1519 -338
rect 1577 -338 1777 -300
rect 1577 -355 1627 -338
rect 1469 -372 1485 -355
rect 1353 -388 1485 -372
rect 1611 -372 1627 -355
rect 1727 -355 1777 -338
rect 1835 -338 2035 -300
rect 1835 -355 1885 -338
rect 1727 -372 1743 -355
rect 1611 -388 1743 -372
rect 1869 -372 1885 -355
rect 1985 -355 2035 -338
rect 2093 -338 2293 -300
rect 2093 -355 2143 -338
rect 1985 -372 2001 -355
rect 1869 -388 2001 -372
rect 2127 -372 2143 -355
rect 2243 -355 2293 -338
rect 2351 -338 2551 -300
rect 2351 -355 2401 -338
rect 2243 -372 2259 -355
rect 2127 -388 2259 -372
rect 2385 -372 2401 -355
rect 2501 -355 2551 -338
rect 2609 -338 2809 -300
rect 2609 -355 2659 -338
rect 2501 -372 2517 -355
rect 2385 -388 2517 -372
rect 2643 -372 2659 -355
rect 2759 -355 2809 -338
rect 2867 -338 3067 -300
rect 2867 -355 2917 -338
rect 2759 -372 2775 -355
rect 2643 -388 2775 -372
rect 2901 -372 2917 -355
rect 3017 -355 3067 -338
rect 3125 -338 3325 -300
rect 3125 -355 3175 -338
rect 3017 -372 3033 -355
rect 2901 -388 3033 -372
rect 3159 -372 3175 -355
rect 3275 -355 3325 -338
rect 3275 -372 3291 -355
rect 3159 -388 3291 -372
<< polycont >>
rect -3275 338 -3175 372
rect -3017 338 -2917 372
rect -2759 338 -2659 372
rect -2501 338 -2401 372
rect -2243 338 -2143 372
rect -1985 338 -1885 372
rect -1727 338 -1627 372
rect -1469 338 -1369 372
rect -1211 338 -1111 372
rect -953 338 -853 372
rect -695 338 -595 372
rect -437 338 -337 372
rect -179 338 -79 372
rect 79 338 179 372
rect 337 338 437 372
rect 595 338 695 372
rect 853 338 953 372
rect 1111 338 1211 372
rect 1369 338 1469 372
rect 1627 338 1727 372
rect 1885 338 1985 372
rect 2143 338 2243 372
rect 2401 338 2501 372
rect 2659 338 2759 372
rect 2917 338 3017 372
rect 3175 338 3275 372
rect -3275 -372 -3175 -338
rect -3017 -372 -2917 -338
rect -2759 -372 -2659 -338
rect -2501 -372 -2401 -338
rect -2243 -372 -2143 -338
rect -1985 -372 -1885 -338
rect -1727 -372 -1627 -338
rect -1469 -372 -1369 -338
rect -1211 -372 -1111 -338
rect -953 -372 -853 -338
rect -695 -372 -595 -338
rect -437 -372 -337 -338
rect -179 -372 -79 -338
rect 79 -372 179 -338
rect 337 -372 437 -338
rect 595 -372 695 -338
rect 853 -372 953 -338
rect 1111 -372 1211 -338
rect 1369 -372 1469 -338
rect 1627 -372 1727 -338
rect 1885 -372 1985 -338
rect 2143 -372 2243 -338
rect 2401 -372 2501 -338
rect 2659 -372 2759 -338
rect 2917 -372 3017 -338
rect 3175 -372 3275 -338
<< locali >>
rect -3505 476 -3409 510
rect 3409 476 3505 510
rect -3505 414 -3471 476
rect 3471 414 3505 476
rect -3291 338 -3275 372
rect -3175 338 -3159 372
rect -3033 338 -3017 372
rect -2917 338 -2901 372
rect -2775 338 -2759 372
rect -2659 338 -2643 372
rect -2517 338 -2501 372
rect -2401 338 -2385 372
rect -2259 338 -2243 372
rect -2143 338 -2127 372
rect -2001 338 -1985 372
rect -1885 338 -1869 372
rect -1743 338 -1727 372
rect -1627 338 -1611 372
rect -1485 338 -1469 372
rect -1369 338 -1353 372
rect -1227 338 -1211 372
rect -1111 338 -1095 372
rect -969 338 -953 372
rect -853 338 -837 372
rect -711 338 -695 372
rect -595 338 -579 372
rect -453 338 -437 372
rect -337 338 -321 372
rect -195 338 -179 372
rect -79 338 -63 372
rect 63 338 79 372
rect 179 338 195 372
rect 321 338 337 372
rect 437 338 453 372
rect 579 338 595 372
rect 695 338 711 372
rect 837 338 853 372
rect 953 338 969 372
rect 1095 338 1111 372
rect 1211 338 1227 372
rect 1353 338 1369 372
rect 1469 338 1485 372
rect 1611 338 1627 372
rect 1727 338 1743 372
rect 1869 338 1885 372
rect 1985 338 2001 372
rect 2127 338 2143 372
rect 2243 338 2259 372
rect 2385 338 2401 372
rect 2501 338 2517 372
rect 2643 338 2659 372
rect 2759 338 2775 372
rect 2901 338 2917 372
rect 3017 338 3033 372
rect 3159 338 3175 372
rect 3275 338 3291 372
rect -3371 288 -3337 304
rect -3371 -304 -3337 -288
rect -3113 288 -3079 304
rect -3113 -304 -3079 -288
rect -2855 288 -2821 304
rect -2855 -304 -2821 -288
rect -2597 288 -2563 304
rect -2597 -304 -2563 -288
rect -2339 288 -2305 304
rect -2339 -304 -2305 -288
rect -2081 288 -2047 304
rect -2081 -304 -2047 -288
rect -1823 288 -1789 304
rect -1823 -304 -1789 -288
rect -1565 288 -1531 304
rect -1565 -304 -1531 -288
rect -1307 288 -1273 304
rect -1307 -304 -1273 -288
rect -1049 288 -1015 304
rect -1049 -304 -1015 -288
rect -791 288 -757 304
rect -791 -304 -757 -288
rect -533 288 -499 304
rect -533 -304 -499 -288
rect -275 288 -241 304
rect -275 -304 -241 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 241 288 275 304
rect 241 -304 275 -288
rect 499 288 533 304
rect 499 -304 533 -288
rect 757 288 791 304
rect 757 -304 791 -288
rect 1015 288 1049 304
rect 1015 -304 1049 -288
rect 1273 288 1307 304
rect 1273 -304 1307 -288
rect 1531 288 1565 304
rect 1531 -304 1565 -288
rect 1789 288 1823 304
rect 1789 -304 1823 -288
rect 2047 288 2081 304
rect 2047 -304 2081 -288
rect 2305 288 2339 304
rect 2305 -304 2339 -288
rect 2563 288 2597 304
rect 2563 -304 2597 -288
rect 2821 288 2855 304
rect 2821 -304 2855 -288
rect 3079 288 3113 304
rect 3079 -304 3113 -288
rect 3337 288 3371 304
rect 3337 -304 3371 -288
rect -3291 -372 -3275 -338
rect -3175 -372 -3159 -338
rect -3033 -372 -3017 -338
rect -2917 -372 -2901 -338
rect -2775 -372 -2759 -338
rect -2659 -372 -2643 -338
rect -2517 -372 -2501 -338
rect -2401 -372 -2385 -338
rect -2259 -372 -2243 -338
rect -2143 -372 -2127 -338
rect -2001 -372 -1985 -338
rect -1885 -372 -1869 -338
rect -1743 -372 -1727 -338
rect -1627 -372 -1611 -338
rect -1485 -372 -1469 -338
rect -1369 -372 -1353 -338
rect -1227 -372 -1211 -338
rect -1111 -372 -1095 -338
rect -969 -372 -953 -338
rect -853 -372 -837 -338
rect -711 -372 -695 -338
rect -595 -372 -579 -338
rect -453 -372 -437 -338
rect -337 -372 -321 -338
rect -195 -372 -179 -338
rect -79 -372 -63 -338
rect 63 -372 79 -338
rect 179 -372 195 -338
rect 321 -372 337 -338
rect 437 -372 453 -338
rect 579 -372 595 -338
rect 695 -372 711 -338
rect 837 -372 853 -338
rect 953 -372 969 -338
rect 1095 -372 1111 -338
rect 1211 -372 1227 -338
rect 1353 -372 1369 -338
rect 1469 -372 1485 -338
rect 1611 -372 1627 -338
rect 1727 -372 1743 -338
rect 1869 -372 1885 -338
rect 1985 -372 2001 -338
rect 2127 -372 2143 -338
rect 2243 -372 2259 -338
rect 2385 -372 2401 -338
rect 2501 -372 2517 -338
rect 2643 -372 2659 -338
rect 2759 -372 2775 -338
rect 2901 -372 2917 -338
rect 3017 -372 3033 -338
rect 3159 -372 3175 -338
rect 3275 -372 3291 -338
rect -3505 -476 -3471 -414
rect 3471 -476 3505 -414
rect -3505 -510 -3409 -476
rect 3409 -510 3505 -476
<< viali >>
rect -3275 338 -3175 372
rect -3017 338 -2917 372
rect -2759 338 -2659 372
rect -2501 338 -2401 372
rect -2243 338 -2143 372
rect -1985 338 -1885 372
rect -1727 338 -1627 372
rect -1469 338 -1369 372
rect -1211 338 -1111 372
rect -953 338 -853 372
rect -695 338 -595 372
rect -437 338 -337 372
rect -179 338 -79 372
rect 79 338 179 372
rect 337 338 437 372
rect 595 338 695 372
rect 853 338 953 372
rect 1111 338 1211 372
rect 1369 338 1469 372
rect 1627 338 1727 372
rect 1885 338 1985 372
rect 2143 338 2243 372
rect 2401 338 2501 372
rect 2659 338 2759 372
rect 2917 338 3017 372
rect 3175 338 3275 372
rect -3371 -288 -3337 288
rect -3113 -288 -3079 288
rect -2855 -288 -2821 288
rect -2597 -288 -2563 288
rect -2339 -288 -2305 288
rect -2081 -288 -2047 288
rect -1823 -288 -1789 288
rect -1565 -288 -1531 288
rect -1307 -288 -1273 288
rect -1049 -288 -1015 288
rect -791 -288 -757 288
rect -533 -288 -499 288
rect -275 -288 -241 288
rect -17 -288 17 288
rect 241 -288 275 288
rect 499 -288 533 288
rect 757 -288 791 288
rect 1015 -288 1049 288
rect 1273 -288 1307 288
rect 1531 -288 1565 288
rect 1789 -288 1823 288
rect 2047 -288 2081 288
rect 2305 -288 2339 288
rect 2563 -288 2597 288
rect 2821 -288 2855 288
rect 3079 -288 3113 288
rect 3337 -288 3371 288
rect -3275 -372 -3175 -338
rect -3017 -372 -2917 -338
rect -2759 -372 -2659 -338
rect -2501 -372 -2401 -338
rect -2243 -372 -2143 -338
rect -1985 -372 -1885 -338
rect -1727 -372 -1627 -338
rect -1469 -372 -1369 -338
rect -1211 -372 -1111 -338
rect -953 -372 -853 -338
rect -695 -372 -595 -338
rect -437 -372 -337 -338
rect -179 -372 -79 -338
rect 79 -372 179 -338
rect 337 -372 437 -338
rect 595 -372 695 -338
rect 853 -372 953 -338
rect 1111 -372 1211 -338
rect 1369 -372 1469 -338
rect 1627 -372 1727 -338
rect 1885 -372 1985 -338
rect 2143 -372 2243 -338
rect 2401 -372 2501 -338
rect 2659 -372 2759 -338
rect 2917 -372 3017 -338
rect 3175 -372 3275 -338
<< metal1 >>
rect -3287 372 -3163 378
rect -3287 338 -3275 372
rect -3175 338 -3163 372
rect -3287 332 -3163 338
rect -3029 372 -2905 378
rect -3029 338 -3017 372
rect -2917 338 -2905 372
rect -3029 332 -2905 338
rect -2771 372 -2647 378
rect -2771 338 -2759 372
rect -2659 338 -2647 372
rect -2771 332 -2647 338
rect -2513 372 -2389 378
rect -2513 338 -2501 372
rect -2401 338 -2389 372
rect -2513 332 -2389 338
rect -2255 372 -2131 378
rect -2255 338 -2243 372
rect -2143 338 -2131 372
rect -2255 332 -2131 338
rect -1997 372 -1873 378
rect -1997 338 -1985 372
rect -1885 338 -1873 372
rect -1997 332 -1873 338
rect -1739 372 -1615 378
rect -1739 338 -1727 372
rect -1627 338 -1615 372
rect -1739 332 -1615 338
rect -1481 372 -1357 378
rect -1481 338 -1469 372
rect -1369 338 -1357 372
rect -1481 332 -1357 338
rect -1223 372 -1099 378
rect -1223 338 -1211 372
rect -1111 338 -1099 372
rect -1223 332 -1099 338
rect -965 372 -841 378
rect -965 338 -953 372
rect -853 338 -841 372
rect -965 332 -841 338
rect -707 372 -583 378
rect -707 338 -695 372
rect -595 338 -583 372
rect -707 332 -583 338
rect -449 372 -325 378
rect -449 338 -437 372
rect -337 338 -325 372
rect -449 332 -325 338
rect -191 372 -67 378
rect -191 338 -179 372
rect -79 338 -67 372
rect -191 332 -67 338
rect 67 372 191 378
rect 67 338 79 372
rect 179 338 191 372
rect 67 332 191 338
rect 325 372 449 378
rect 325 338 337 372
rect 437 338 449 372
rect 325 332 449 338
rect 583 372 707 378
rect 583 338 595 372
rect 695 338 707 372
rect 583 332 707 338
rect 841 372 965 378
rect 841 338 853 372
rect 953 338 965 372
rect 841 332 965 338
rect 1099 372 1223 378
rect 1099 338 1111 372
rect 1211 338 1223 372
rect 1099 332 1223 338
rect 1357 372 1481 378
rect 1357 338 1369 372
rect 1469 338 1481 372
rect 1357 332 1481 338
rect 1615 372 1739 378
rect 1615 338 1627 372
rect 1727 338 1739 372
rect 1615 332 1739 338
rect 1873 372 1997 378
rect 1873 338 1885 372
rect 1985 338 1997 372
rect 1873 332 1997 338
rect 2131 372 2255 378
rect 2131 338 2143 372
rect 2243 338 2255 372
rect 2131 332 2255 338
rect 2389 372 2513 378
rect 2389 338 2401 372
rect 2501 338 2513 372
rect 2389 332 2513 338
rect 2647 372 2771 378
rect 2647 338 2659 372
rect 2759 338 2771 372
rect 2647 332 2771 338
rect 2905 372 3029 378
rect 2905 338 2917 372
rect 3017 338 3029 372
rect 2905 332 3029 338
rect 3163 372 3287 378
rect 3163 338 3175 372
rect 3275 338 3287 372
rect 3163 332 3287 338
rect -3377 288 -3331 300
rect -3377 -288 -3371 288
rect -3337 -288 -3331 288
rect -3377 -300 -3331 -288
rect -3119 288 -3073 300
rect -3119 -288 -3113 288
rect -3079 -288 -3073 288
rect -3119 -300 -3073 -288
rect -2861 288 -2815 300
rect -2861 -288 -2855 288
rect -2821 -288 -2815 288
rect -2861 -300 -2815 -288
rect -2603 288 -2557 300
rect -2603 -288 -2597 288
rect -2563 -288 -2557 288
rect -2603 -300 -2557 -288
rect -2345 288 -2299 300
rect -2345 -288 -2339 288
rect -2305 -288 -2299 288
rect -2345 -300 -2299 -288
rect -2087 288 -2041 300
rect -2087 -288 -2081 288
rect -2047 -288 -2041 288
rect -2087 -300 -2041 -288
rect -1829 288 -1783 300
rect -1829 -288 -1823 288
rect -1789 -288 -1783 288
rect -1829 -300 -1783 -288
rect -1571 288 -1525 300
rect -1571 -288 -1565 288
rect -1531 -288 -1525 288
rect -1571 -300 -1525 -288
rect -1313 288 -1267 300
rect -1313 -288 -1307 288
rect -1273 -288 -1267 288
rect -1313 -300 -1267 -288
rect -1055 288 -1009 300
rect -1055 -288 -1049 288
rect -1015 -288 -1009 288
rect -1055 -300 -1009 -288
rect -797 288 -751 300
rect -797 -288 -791 288
rect -757 -288 -751 288
rect -797 -300 -751 -288
rect -539 288 -493 300
rect -539 -288 -533 288
rect -499 -288 -493 288
rect -539 -300 -493 -288
rect -281 288 -235 300
rect -281 -288 -275 288
rect -241 -288 -235 288
rect -281 -300 -235 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 235 288 281 300
rect 235 -288 241 288
rect 275 -288 281 288
rect 235 -300 281 -288
rect 493 288 539 300
rect 493 -288 499 288
rect 533 -288 539 288
rect 493 -300 539 -288
rect 751 288 797 300
rect 751 -288 757 288
rect 791 -288 797 288
rect 751 -300 797 -288
rect 1009 288 1055 300
rect 1009 -288 1015 288
rect 1049 -288 1055 288
rect 1009 -300 1055 -288
rect 1267 288 1313 300
rect 1267 -288 1273 288
rect 1307 -288 1313 288
rect 1267 -300 1313 -288
rect 1525 288 1571 300
rect 1525 -288 1531 288
rect 1565 -288 1571 288
rect 1525 -300 1571 -288
rect 1783 288 1829 300
rect 1783 -288 1789 288
rect 1823 -288 1829 288
rect 1783 -300 1829 -288
rect 2041 288 2087 300
rect 2041 -288 2047 288
rect 2081 -288 2087 288
rect 2041 -300 2087 -288
rect 2299 288 2345 300
rect 2299 -288 2305 288
rect 2339 -288 2345 288
rect 2299 -300 2345 -288
rect 2557 288 2603 300
rect 2557 -288 2563 288
rect 2597 -288 2603 288
rect 2557 -300 2603 -288
rect 2815 288 2861 300
rect 2815 -288 2821 288
rect 2855 -288 2861 288
rect 2815 -300 2861 -288
rect 3073 288 3119 300
rect 3073 -288 3079 288
rect 3113 -288 3119 288
rect 3073 -300 3119 -288
rect 3331 288 3377 300
rect 3331 -288 3337 288
rect 3371 -288 3377 288
rect 3331 -300 3377 -288
rect -3287 -338 -3163 -332
rect -3287 -372 -3275 -338
rect -3175 -372 -3163 -338
rect -3287 -378 -3163 -372
rect -3029 -338 -2905 -332
rect -3029 -372 -3017 -338
rect -2917 -372 -2905 -338
rect -3029 -378 -2905 -372
rect -2771 -338 -2647 -332
rect -2771 -372 -2759 -338
rect -2659 -372 -2647 -338
rect -2771 -378 -2647 -372
rect -2513 -338 -2389 -332
rect -2513 -372 -2501 -338
rect -2401 -372 -2389 -338
rect -2513 -378 -2389 -372
rect -2255 -338 -2131 -332
rect -2255 -372 -2243 -338
rect -2143 -372 -2131 -338
rect -2255 -378 -2131 -372
rect -1997 -338 -1873 -332
rect -1997 -372 -1985 -338
rect -1885 -372 -1873 -338
rect -1997 -378 -1873 -372
rect -1739 -338 -1615 -332
rect -1739 -372 -1727 -338
rect -1627 -372 -1615 -338
rect -1739 -378 -1615 -372
rect -1481 -338 -1357 -332
rect -1481 -372 -1469 -338
rect -1369 -372 -1357 -338
rect -1481 -378 -1357 -372
rect -1223 -338 -1099 -332
rect -1223 -372 -1211 -338
rect -1111 -372 -1099 -338
rect -1223 -378 -1099 -372
rect -965 -338 -841 -332
rect -965 -372 -953 -338
rect -853 -372 -841 -338
rect -965 -378 -841 -372
rect -707 -338 -583 -332
rect -707 -372 -695 -338
rect -595 -372 -583 -338
rect -707 -378 -583 -372
rect -449 -338 -325 -332
rect -449 -372 -437 -338
rect -337 -372 -325 -338
rect -449 -378 -325 -372
rect -191 -338 -67 -332
rect -191 -372 -179 -338
rect -79 -372 -67 -338
rect -191 -378 -67 -372
rect 67 -338 191 -332
rect 67 -372 79 -338
rect 179 -372 191 -338
rect 67 -378 191 -372
rect 325 -338 449 -332
rect 325 -372 337 -338
rect 437 -372 449 -338
rect 325 -378 449 -372
rect 583 -338 707 -332
rect 583 -372 595 -338
rect 695 -372 707 -338
rect 583 -378 707 -372
rect 841 -338 965 -332
rect 841 -372 853 -338
rect 953 -372 965 -338
rect 841 -378 965 -372
rect 1099 -338 1223 -332
rect 1099 -372 1111 -338
rect 1211 -372 1223 -338
rect 1099 -378 1223 -372
rect 1357 -338 1481 -332
rect 1357 -372 1369 -338
rect 1469 -372 1481 -338
rect 1357 -378 1481 -372
rect 1615 -338 1739 -332
rect 1615 -372 1627 -338
rect 1727 -372 1739 -338
rect 1615 -378 1739 -372
rect 1873 -338 1997 -332
rect 1873 -372 1885 -338
rect 1985 -372 1997 -338
rect 1873 -378 1997 -372
rect 2131 -338 2255 -332
rect 2131 -372 2143 -338
rect 2243 -372 2255 -338
rect 2131 -378 2255 -372
rect 2389 -338 2513 -332
rect 2389 -372 2401 -338
rect 2501 -372 2513 -338
rect 2389 -378 2513 -372
rect 2647 -338 2771 -332
rect 2647 -372 2659 -338
rect 2759 -372 2771 -338
rect 2647 -378 2771 -372
rect 2905 -338 3029 -332
rect 2905 -372 2917 -338
rect 3017 -372 3029 -338
rect 2905 -378 3029 -372
rect 3163 -338 3287 -332
rect 3163 -372 3175 -338
rect 3275 -372 3287 -338
rect 3163 -378 3287 -372
<< properties >>
string FIXED_BBOX -3488 -493 3488 493
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3 l 1 m 1 nf 26 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713300419
<< pwell >>
rect -3553 -858 3553 858
<< mvnmos >>
rect -3325 -600 -3125 600
rect -3067 -600 -2867 600
rect -2809 -600 -2609 600
rect -2551 -600 -2351 600
rect -2293 -600 -2093 600
rect -2035 -600 -1835 600
rect -1777 -600 -1577 600
rect -1519 -600 -1319 600
rect -1261 -600 -1061 600
rect -1003 -600 -803 600
rect -745 -600 -545 600
rect -487 -600 -287 600
rect -229 -600 -29 600
rect 29 -600 229 600
rect 287 -600 487 600
rect 545 -600 745 600
rect 803 -600 1003 600
rect 1061 -600 1261 600
rect 1319 -600 1519 600
rect 1577 -600 1777 600
rect 1835 -600 2035 600
rect 2093 -600 2293 600
rect 2351 -600 2551 600
rect 2609 -600 2809 600
rect 2867 -600 3067 600
rect 3125 -600 3325 600
<< mvndiff >>
rect -3383 588 -3325 600
rect -3383 -588 -3371 588
rect -3337 -588 -3325 588
rect -3383 -600 -3325 -588
rect -3125 588 -3067 600
rect -3125 -588 -3113 588
rect -3079 -588 -3067 588
rect -3125 -600 -3067 -588
rect -2867 588 -2809 600
rect -2867 -588 -2855 588
rect -2821 -588 -2809 588
rect -2867 -600 -2809 -588
rect -2609 588 -2551 600
rect -2609 -588 -2597 588
rect -2563 -588 -2551 588
rect -2609 -600 -2551 -588
rect -2351 588 -2293 600
rect -2351 -588 -2339 588
rect -2305 -588 -2293 588
rect -2351 -600 -2293 -588
rect -2093 588 -2035 600
rect -2093 -588 -2081 588
rect -2047 -588 -2035 588
rect -2093 -600 -2035 -588
rect -1835 588 -1777 600
rect -1835 -588 -1823 588
rect -1789 -588 -1777 588
rect -1835 -600 -1777 -588
rect -1577 588 -1519 600
rect -1577 -588 -1565 588
rect -1531 -588 -1519 588
rect -1577 -600 -1519 -588
rect -1319 588 -1261 600
rect -1319 -588 -1307 588
rect -1273 -588 -1261 588
rect -1319 -600 -1261 -588
rect -1061 588 -1003 600
rect -1061 -588 -1049 588
rect -1015 -588 -1003 588
rect -1061 -600 -1003 -588
rect -803 588 -745 600
rect -803 -588 -791 588
rect -757 -588 -745 588
rect -803 -600 -745 -588
rect -545 588 -487 600
rect -545 -588 -533 588
rect -499 -588 -487 588
rect -545 -600 -487 -588
rect -287 588 -229 600
rect -287 -588 -275 588
rect -241 -588 -229 588
rect -287 -600 -229 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 229 588 287 600
rect 229 -588 241 588
rect 275 -588 287 588
rect 229 -600 287 -588
rect 487 588 545 600
rect 487 -588 499 588
rect 533 -588 545 588
rect 487 -600 545 -588
rect 745 588 803 600
rect 745 -588 757 588
rect 791 -588 803 588
rect 745 -600 803 -588
rect 1003 588 1061 600
rect 1003 -588 1015 588
rect 1049 -588 1061 588
rect 1003 -600 1061 -588
rect 1261 588 1319 600
rect 1261 -588 1273 588
rect 1307 -588 1319 588
rect 1261 -600 1319 -588
rect 1519 588 1577 600
rect 1519 -588 1531 588
rect 1565 -588 1577 588
rect 1519 -600 1577 -588
rect 1777 588 1835 600
rect 1777 -588 1789 588
rect 1823 -588 1835 588
rect 1777 -600 1835 -588
rect 2035 588 2093 600
rect 2035 -588 2047 588
rect 2081 -588 2093 588
rect 2035 -600 2093 -588
rect 2293 588 2351 600
rect 2293 -588 2305 588
rect 2339 -588 2351 588
rect 2293 -600 2351 -588
rect 2551 588 2609 600
rect 2551 -588 2563 588
rect 2597 -588 2609 588
rect 2551 -600 2609 -588
rect 2809 588 2867 600
rect 2809 -588 2821 588
rect 2855 -588 2867 588
rect 2809 -600 2867 -588
rect 3067 588 3125 600
rect 3067 -588 3079 588
rect 3113 -588 3125 588
rect 3067 -600 3125 -588
rect 3325 588 3383 600
rect 3325 -588 3337 588
rect 3371 -588 3383 588
rect 3325 -600 3383 -588
<< mvndiffc >>
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
<< mvpsubdiff >>
rect -3517 810 3517 822
rect -3517 776 -3409 810
rect 3409 776 3517 810
rect -3517 764 3517 776
rect -3517 714 -3459 764
rect -3517 -714 -3505 714
rect -3471 -714 -3459 714
rect 3459 714 3517 764
rect -3517 -764 -3459 -714
rect 3459 -714 3471 714
rect 3505 -714 3517 714
rect 3459 -764 3517 -714
rect -3517 -776 3517 -764
rect -3517 -810 -3409 -776
rect 3409 -810 3517 -776
rect -3517 -822 3517 -810
<< mvpsubdiffcont >>
rect -3409 776 3409 810
rect -3505 -714 -3471 714
rect 3471 -714 3505 714
rect -3409 -810 3409 -776
<< poly >>
rect -3291 672 -3159 688
rect -3291 655 -3275 672
rect -3325 638 -3275 655
rect -3175 655 -3159 672
rect -3033 672 -2901 688
rect -3033 655 -3017 672
rect -3175 638 -3125 655
rect -3325 600 -3125 638
rect -3067 638 -3017 655
rect -2917 655 -2901 672
rect -2775 672 -2643 688
rect -2775 655 -2759 672
rect -2917 638 -2867 655
rect -3067 600 -2867 638
rect -2809 638 -2759 655
rect -2659 655 -2643 672
rect -2517 672 -2385 688
rect -2517 655 -2501 672
rect -2659 638 -2609 655
rect -2809 600 -2609 638
rect -2551 638 -2501 655
rect -2401 655 -2385 672
rect -2259 672 -2127 688
rect -2259 655 -2243 672
rect -2401 638 -2351 655
rect -2551 600 -2351 638
rect -2293 638 -2243 655
rect -2143 655 -2127 672
rect -2001 672 -1869 688
rect -2001 655 -1985 672
rect -2143 638 -2093 655
rect -2293 600 -2093 638
rect -2035 638 -1985 655
rect -1885 655 -1869 672
rect -1743 672 -1611 688
rect -1743 655 -1727 672
rect -1885 638 -1835 655
rect -2035 600 -1835 638
rect -1777 638 -1727 655
rect -1627 655 -1611 672
rect -1485 672 -1353 688
rect -1485 655 -1469 672
rect -1627 638 -1577 655
rect -1777 600 -1577 638
rect -1519 638 -1469 655
rect -1369 655 -1353 672
rect -1227 672 -1095 688
rect -1227 655 -1211 672
rect -1369 638 -1319 655
rect -1519 600 -1319 638
rect -1261 638 -1211 655
rect -1111 655 -1095 672
rect -969 672 -837 688
rect -969 655 -953 672
rect -1111 638 -1061 655
rect -1261 600 -1061 638
rect -1003 638 -953 655
rect -853 655 -837 672
rect -711 672 -579 688
rect -711 655 -695 672
rect -853 638 -803 655
rect -1003 600 -803 638
rect -745 638 -695 655
rect -595 655 -579 672
rect -453 672 -321 688
rect -453 655 -437 672
rect -595 638 -545 655
rect -745 600 -545 638
rect -487 638 -437 655
rect -337 655 -321 672
rect -195 672 -63 688
rect -195 655 -179 672
rect -337 638 -287 655
rect -487 600 -287 638
rect -229 638 -179 655
rect -79 655 -63 672
rect 63 672 195 688
rect 63 655 79 672
rect -79 638 -29 655
rect -229 600 -29 638
rect 29 638 79 655
rect 179 655 195 672
rect 321 672 453 688
rect 321 655 337 672
rect 179 638 229 655
rect 29 600 229 638
rect 287 638 337 655
rect 437 655 453 672
rect 579 672 711 688
rect 579 655 595 672
rect 437 638 487 655
rect 287 600 487 638
rect 545 638 595 655
rect 695 655 711 672
rect 837 672 969 688
rect 837 655 853 672
rect 695 638 745 655
rect 545 600 745 638
rect 803 638 853 655
rect 953 655 969 672
rect 1095 672 1227 688
rect 1095 655 1111 672
rect 953 638 1003 655
rect 803 600 1003 638
rect 1061 638 1111 655
rect 1211 655 1227 672
rect 1353 672 1485 688
rect 1353 655 1369 672
rect 1211 638 1261 655
rect 1061 600 1261 638
rect 1319 638 1369 655
rect 1469 655 1485 672
rect 1611 672 1743 688
rect 1611 655 1627 672
rect 1469 638 1519 655
rect 1319 600 1519 638
rect 1577 638 1627 655
rect 1727 655 1743 672
rect 1869 672 2001 688
rect 1869 655 1885 672
rect 1727 638 1777 655
rect 1577 600 1777 638
rect 1835 638 1885 655
rect 1985 655 2001 672
rect 2127 672 2259 688
rect 2127 655 2143 672
rect 1985 638 2035 655
rect 1835 600 2035 638
rect 2093 638 2143 655
rect 2243 655 2259 672
rect 2385 672 2517 688
rect 2385 655 2401 672
rect 2243 638 2293 655
rect 2093 600 2293 638
rect 2351 638 2401 655
rect 2501 655 2517 672
rect 2643 672 2775 688
rect 2643 655 2659 672
rect 2501 638 2551 655
rect 2351 600 2551 638
rect 2609 638 2659 655
rect 2759 655 2775 672
rect 2901 672 3033 688
rect 2901 655 2917 672
rect 2759 638 2809 655
rect 2609 600 2809 638
rect 2867 638 2917 655
rect 3017 655 3033 672
rect 3159 672 3291 688
rect 3159 655 3175 672
rect 3017 638 3067 655
rect 2867 600 3067 638
rect 3125 638 3175 655
rect 3275 655 3291 672
rect 3275 638 3325 655
rect 3125 600 3325 638
rect -3325 -638 -3125 -600
rect -3325 -655 -3275 -638
rect -3291 -672 -3275 -655
rect -3175 -655 -3125 -638
rect -3067 -638 -2867 -600
rect -3067 -655 -3017 -638
rect -3175 -672 -3159 -655
rect -3291 -688 -3159 -672
rect -3033 -672 -3017 -655
rect -2917 -655 -2867 -638
rect -2809 -638 -2609 -600
rect -2809 -655 -2759 -638
rect -2917 -672 -2901 -655
rect -3033 -688 -2901 -672
rect -2775 -672 -2759 -655
rect -2659 -655 -2609 -638
rect -2551 -638 -2351 -600
rect -2551 -655 -2501 -638
rect -2659 -672 -2643 -655
rect -2775 -688 -2643 -672
rect -2517 -672 -2501 -655
rect -2401 -655 -2351 -638
rect -2293 -638 -2093 -600
rect -2293 -655 -2243 -638
rect -2401 -672 -2385 -655
rect -2517 -688 -2385 -672
rect -2259 -672 -2243 -655
rect -2143 -655 -2093 -638
rect -2035 -638 -1835 -600
rect -2035 -655 -1985 -638
rect -2143 -672 -2127 -655
rect -2259 -688 -2127 -672
rect -2001 -672 -1985 -655
rect -1885 -655 -1835 -638
rect -1777 -638 -1577 -600
rect -1777 -655 -1727 -638
rect -1885 -672 -1869 -655
rect -2001 -688 -1869 -672
rect -1743 -672 -1727 -655
rect -1627 -655 -1577 -638
rect -1519 -638 -1319 -600
rect -1519 -655 -1469 -638
rect -1627 -672 -1611 -655
rect -1743 -688 -1611 -672
rect -1485 -672 -1469 -655
rect -1369 -655 -1319 -638
rect -1261 -638 -1061 -600
rect -1261 -655 -1211 -638
rect -1369 -672 -1353 -655
rect -1485 -688 -1353 -672
rect -1227 -672 -1211 -655
rect -1111 -655 -1061 -638
rect -1003 -638 -803 -600
rect -1003 -655 -953 -638
rect -1111 -672 -1095 -655
rect -1227 -688 -1095 -672
rect -969 -672 -953 -655
rect -853 -655 -803 -638
rect -745 -638 -545 -600
rect -745 -655 -695 -638
rect -853 -672 -837 -655
rect -969 -688 -837 -672
rect -711 -672 -695 -655
rect -595 -655 -545 -638
rect -487 -638 -287 -600
rect -487 -655 -437 -638
rect -595 -672 -579 -655
rect -711 -688 -579 -672
rect -453 -672 -437 -655
rect -337 -655 -287 -638
rect -229 -638 -29 -600
rect -229 -655 -179 -638
rect -337 -672 -321 -655
rect -453 -688 -321 -672
rect -195 -672 -179 -655
rect -79 -655 -29 -638
rect 29 -638 229 -600
rect 29 -655 79 -638
rect -79 -672 -63 -655
rect -195 -688 -63 -672
rect 63 -672 79 -655
rect 179 -655 229 -638
rect 287 -638 487 -600
rect 287 -655 337 -638
rect 179 -672 195 -655
rect 63 -688 195 -672
rect 321 -672 337 -655
rect 437 -655 487 -638
rect 545 -638 745 -600
rect 545 -655 595 -638
rect 437 -672 453 -655
rect 321 -688 453 -672
rect 579 -672 595 -655
rect 695 -655 745 -638
rect 803 -638 1003 -600
rect 803 -655 853 -638
rect 695 -672 711 -655
rect 579 -688 711 -672
rect 837 -672 853 -655
rect 953 -655 1003 -638
rect 1061 -638 1261 -600
rect 1061 -655 1111 -638
rect 953 -672 969 -655
rect 837 -688 969 -672
rect 1095 -672 1111 -655
rect 1211 -655 1261 -638
rect 1319 -638 1519 -600
rect 1319 -655 1369 -638
rect 1211 -672 1227 -655
rect 1095 -688 1227 -672
rect 1353 -672 1369 -655
rect 1469 -655 1519 -638
rect 1577 -638 1777 -600
rect 1577 -655 1627 -638
rect 1469 -672 1485 -655
rect 1353 -688 1485 -672
rect 1611 -672 1627 -655
rect 1727 -655 1777 -638
rect 1835 -638 2035 -600
rect 1835 -655 1885 -638
rect 1727 -672 1743 -655
rect 1611 -688 1743 -672
rect 1869 -672 1885 -655
rect 1985 -655 2035 -638
rect 2093 -638 2293 -600
rect 2093 -655 2143 -638
rect 1985 -672 2001 -655
rect 1869 -688 2001 -672
rect 2127 -672 2143 -655
rect 2243 -655 2293 -638
rect 2351 -638 2551 -600
rect 2351 -655 2401 -638
rect 2243 -672 2259 -655
rect 2127 -688 2259 -672
rect 2385 -672 2401 -655
rect 2501 -655 2551 -638
rect 2609 -638 2809 -600
rect 2609 -655 2659 -638
rect 2501 -672 2517 -655
rect 2385 -688 2517 -672
rect 2643 -672 2659 -655
rect 2759 -655 2809 -638
rect 2867 -638 3067 -600
rect 2867 -655 2917 -638
rect 2759 -672 2775 -655
rect 2643 -688 2775 -672
rect 2901 -672 2917 -655
rect 3017 -655 3067 -638
rect 3125 -638 3325 -600
rect 3125 -655 3175 -638
rect 3017 -672 3033 -655
rect 2901 -688 3033 -672
rect 3159 -672 3175 -655
rect 3275 -655 3325 -638
rect 3275 -672 3291 -655
rect 3159 -688 3291 -672
<< polycont >>
rect -3275 638 -3175 672
rect -3017 638 -2917 672
rect -2759 638 -2659 672
rect -2501 638 -2401 672
rect -2243 638 -2143 672
rect -1985 638 -1885 672
rect -1727 638 -1627 672
rect -1469 638 -1369 672
rect -1211 638 -1111 672
rect -953 638 -853 672
rect -695 638 -595 672
rect -437 638 -337 672
rect -179 638 -79 672
rect 79 638 179 672
rect 337 638 437 672
rect 595 638 695 672
rect 853 638 953 672
rect 1111 638 1211 672
rect 1369 638 1469 672
rect 1627 638 1727 672
rect 1885 638 1985 672
rect 2143 638 2243 672
rect 2401 638 2501 672
rect 2659 638 2759 672
rect 2917 638 3017 672
rect 3175 638 3275 672
rect -3275 -672 -3175 -638
rect -3017 -672 -2917 -638
rect -2759 -672 -2659 -638
rect -2501 -672 -2401 -638
rect -2243 -672 -2143 -638
rect -1985 -672 -1885 -638
rect -1727 -672 -1627 -638
rect -1469 -672 -1369 -638
rect -1211 -672 -1111 -638
rect -953 -672 -853 -638
rect -695 -672 -595 -638
rect -437 -672 -337 -638
rect -179 -672 -79 -638
rect 79 -672 179 -638
rect 337 -672 437 -638
rect 595 -672 695 -638
rect 853 -672 953 -638
rect 1111 -672 1211 -638
rect 1369 -672 1469 -638
rect 1627 -672 1727 -638
rect 1885 -672 1985 -638
rect 2143 -672 2243 -638
rect 2401 -672 2501 -638
rect 2659 -672 2759 -638
rect 2917 -672 3017 -638
rect 3175 -672 3275 -638
<< locali >>
rect -3505 776 -3409 810
rect 3409 776 3505 810
rect -3505 714 -3471 776
rect 3471 714 3505 776
rect -3291 638 -3275 672
rect -3175 638 -3159 672
rect -3033 638 -3017 672
rect -2917 638 -2901 672
rect -2775 638 -2759 672
rect -2659 638 -2643 672
rect -2517 638 -2501 672
rect -2401 638 -2385 672
rect -2259 638 -2243 672
rect -2143 638 -2127 672
rect -2001 638 -1985 672
rect -1885 638 -1869 672
rect -1743 638 -1727 672
rect -1627 638 -1611 672
rect -1485 638 -1469 672
rect -1369 638 -1353 672
rect -1227 638 -1211 672
rect -1111 638 -1095 672
rect -969 638 -953 672
rect -853 638 -837 672
rect -711 638 -695 672
rect -595 638 -579 672
rect -453 638 -437 672
rect -337 638 -321 672
rect -195 638 -179 672
rect -79 638 -63 672
rect 63 638 79 672
rect 179 638 195 672
rect 321 638 337 672
rect 437 638 453 672
rect 579 638 595 672
rect 695 638 711 672
rect 837 638 853 672
rect 953 638 969 672
rect 1095 638 1111 672
rect 1211 638 1227 672
rect 1353 638 1369 672
rect 1469 638 1485 672
rect 1611 638 1627 672
rect 1727 638 1743 672
rect 1869 638 1885 672
rect 1985 638 2001 672
rect 2127 638 2143 672
rect 2243 638 2259 672
rect 2385 638 2401 672
rect 2501 638 2517 672
rect 2643 638 2659 672
rect 2759 638 2775 672
rect 2901 638 2917 672
rect 3017 638 3033 672
rect 3159 638 3175 672
rect 3275 638 3291 672
rect -3371 588 -3337 604
rect -3371 -604 -3337 -588
rect -3113 588 -3079 604
rect -3113 -604 -3079 -588
rect -2855 588 -2821 604
rect -2855 -604 -2821 -588
rect -2597 588 -2563 604
rect -2597 -604 -2563 -588
rect -2339 588 -2305 604
rect -2339 -604 -2305 -588
rect -2081 588 -2047 604
rect -2081 -604 -2047 -588
rect -1823 588 -1789 604
rect -1823 -604 -1789 -588
rect -1565 588 -1531 604
rect -1565 -604 -1531 -588
rect -1307 588 -1273 604
rect -1307 -604 -1273 -588
rect -1049 588 -1015 604
rect -1049 -604 -1015 -588
rect -791 588 -757 604
rect -791 -604 -757 -588
rect -533 588 -499 604
rect -533 -604 -499 -588
rect -275 588 -241 604
rect -275 -604 -241 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 241 588 275 604
rect 241 -604 275 -588
rect 499 588 533 604
rect 499 -604 533 -588
rect 757 588 791 604
rect 757 -604 791 -588
rect 1015 588 1049 604
rect 1015 -604 1049 -588
rect 1273 588 1307 604
rect 1273 -604 1307 -588
rect 1531 588 1565 604
rect 1531 -604 1565 -588
rect 1789 588 1823 604
rect 1789 -604 1823 -588
rect 2047 588 2081 604
rect 2047 -604 2081 -588
rect 2305 588 2339 604
rect 2305 -604 2339 -588
rect 2563 588 2597 604
rect 2563 -604 2597 -588
rect 2821 588 2855 604
rect 2821 -604 2855 -588
rect 3079 588 3113 604
rect 3079 -604 3113 -588
rect 3337 588 3371 604
rect 3337 -604 3371 -588
rect -3291 -672 -3275 -638
rect -3175 -672 -3159 -638
rect -3033 -672 -3017 -638
rect -2917 -672 -2901 -638
rect -2775 -672 -2759 -638
rect -2659 -672 -2643 -638
rect -2517 -672 -2501 -638
rect -2401 -672 -2385 -638
rect -2259 -672 -2243 -638
rect -2143 -672 -2127 -638
rect -2001 -672 -1985 -638
rect -1885 -672 -1869 -638
rect -1743 -672 -1727 -638
rect -1627 -672 -1611 -638
rect -1485 -672 -1469 -638
rect -1369 -672 -1353 -638
rect -1227 -672 -1211 -638
rect -1111 -672 -1095 -638
rect -969 -672 -953 -638
rect -853 -672 -837 -638
rect -711 -672 -695 -638
rect -595 -672 -579 -638
rect -453 -672 -437 -638
rect -337 -672 -321 -638
rect -195 -672 -179 -638
rect -79 -672 -63 -638
rect 63 -672 79 -638
rect 179 -672 195 -638
rect 321 -672 337 -638
rect 437 -672 453 -638
rect 579 -672 595 -638
rect 695 -672 711 -638
rect 837 -672 853 -638
rect 953 -672 969 -638
rect 1095 -672 1111 -638
rect 1211 -672 1227 -638
rect 1353 -672 1369 -638
rect 1469 -672 1485 -638
rect 1611 -672 1627 -638
rect 1727 -672 1743 -638
rect 1869 -672 1885 -638
rect 1985 -672 2001 -638
rect 2127 -672 2143 -638
rect 2243 -672 2259 -638
rect 2385 -672 2401 -638
rect 2501 -672 2517 -638
rect 2643 -672 2659 -638
rect 2759 -672 2775 -638
rect 2901 -672 2917 -638
rect 3017 -672 3033 -638
rect 3159 -672 3175 -638
rect 3275 -672 3291 -638
rect -3505 -776 -3471 -714
rect 3471 -776 3505 -714
rect -3505 -810 -3409 -776
rect 3409 -810 3505 -776
<< viali >>
rect -3275 638 -3175 672
rect -3017 638 -2917 672
rect -2759 638 -2659 672
rect -2501 638 -2401 672
rect -2243 638 -2143 672
rect -1985 638 -1885 672
rect -1727 638 -1627 672
rect -1469 638 -1369 672
rect -1211 638 -1111 672
rect -953 638 -853 672
rect -695 638 -595 672
rect -437 638 -337 672
rect -179 638 -79 672
rect 79 638 179 672
rect 337 638 437 672
rect 595 638 695 672
rect 853 638 953 672
rect 1111 638 1211 672
rect 1369 638 1469 672
rect 1627 638 1727 672
rect 1885 638 1985 672
rect 2143 638 2243 672
rect 2401 638 2501 672
rect 2659 638 2759 672
rect 2917 638 3017 672
rect 3175 638 3275 672
rect -3371 -588 -3337 588
rect -3113 -588 -3079 588
rect -2855 -588 -2821 588
rect -2597 -588 -2563 588
rect -2339 -588 -2305 588
rect -2081 -588 -2047 588
rect -1823 -588 -1789 588
rect -1565 -588 -1531 588
rect -1307 -588 -1273 588
rect -1049 -588 -1015 588
rect -791 -588 -757 588
rect -533 -588 -499 588
rect -275 -588 -241 588
rect -17 -588 17 588
rect 241 -588 275 588
rect 499 -588 533 588
rect 757 -588 791 588
rect 1015 -588 1049 588
rect 1273 -588 1307 588
rect 1531 -588 1565 588
rect 1789 -588 1823 588
rect 2047 -588 2081 588
rect 2305 -588 2339 588
rect 2563 -588 2597 588
rect 2821 -588 2855 588
rect 3079 -588 3113 588
rect 3337 -588 3371 588
rect -3275 -672 -3175 -638
rect -3017 -672 -2917 -638
rect -2759 -672 -2659 -638
rect -2501 -672 -2401 -638
rect -2243 -672 -2143 -638
rect -1985 -672 -1885 -638
rect -1727 -672 -1627 -638
rect -1469 -672 -1369 -638
rect -1211 -672 -1111 -638
rect -953 -672 -853 -638
rect -695 -672 -595 -638
rect -437 -672 -337 -638
rect -179 -672 -79 -638
rect 79 -672 179 -638
rect 337 -672 437 -638
rect 595 -672 695 -638
rect 853 -672 953 -638
rect 1111 -672 1211 -638
rect 1369 -672 1469 -638
rect 1627 -672 1727 -638
rect 1885 -672 1985 -638
rect 2143 -672 2243 -638
rect 2401 -672 2501 -638
rect 2659 -672 2759 -638
rect 2917 -672 3017 -638
rect 3175 -672 3275 -638
<< metal1 >>
rect -3287 672 -3163 678
rect -3287 638 -3275 672
rect -3175 638 -3163 672
rect -3287 632 -3163 638
rect -3029 672 -2905 678
rect -3029 638 -3017 672
rect -2917 638 -2905 672
rect -3029 632 -2905 638
rect -2771 672 -2647 678
rect -2771 638 -2759 672
rect -2659 638 -2647 672
rect -2771 632 -2647 638
rect -2513 672 -2389 678
rect -2513 638 -2501 672
rect -2401 638 -2389 672
rect -2513 632 -2389 638
rect -2255 672 -2131 678
rect -2255 638 -2243 672
rect -2143 638 -2131 672
rect -2255 632 -2131 638
rect -1997 672 -1873 678
rect -1997 638 -1985 672
rect -1885 638 -1873 672
rect -1997 632 -1873 638
rect -1739 672 -1615 678
rect -1739 638 -1727 672
rect -1627 638 -1615 672
rect -1739 632 -1615 638
rect -1481 672 -1357 678
rect -1481 638 -1469 672
rect -1369 638 -1357 672
rect -1481 632 -1357 638
rect -1223 672 -1099 678
rect -1223 638 -1211 672
rect -1111 638 -1099 672
rect -1223 632 -1099 638
rect -965 672 -841 678
rect -965 638 -953 672
rect -853 638 -841 672
rect -965 632 -841 638
rect -707 672 -583 678
rect -707 638 -695 672
rect -595 638 -583 672
rect -707 632 -583 638
rect -449 672 -325 678
rect -449 638 -437 672
rect -337 638 -325 672
rect -449 632 -325 638
rect -191 672 -67 678
rect -191 638 -179 672
rect -79 638 -67 672
rect -191 632 -67 638
rect 67 672 191 678
rect 67 638 79 672
rect 179 638 191 672
rect 67 632 191 638
rect 325 672 449 678
rect 325 638 337 672
rect 437 638 449 672
rect 325 632 449 638
rect 583 672 707 678
rect 583 638 595 672
rect 695 638 707 672
rect 583 632 707 638
rect 841 672 965 678
rect 841 638 853 672
rect 953 638 965 672
rect 841 632 965 638
rect 1099 672 1223 678
rect 1099 638 1111 672
rect 1211 638 1223 672
rect 1099 632 1223 638
rect 1357 672 1481 678
rect 1357 638 1369 672
rect 1469 638 1481 672
rect 1357 632 1481 638
rect 1615 672 1739 678
rect 1615 638 1627 672
rect 1727 638 1739 672
rect 1615 632 1739 638
rect 1873 672 1997 678
rect 1873 638 1885 672
rect 1985 638 1997 672
rect 1873 632 1997 638
rect 2131 672 2255 678
rect 2131 638 2143 672
rect 2243 638 2255 672
rect 2131 632 2255 638
rect 2389 672 2513 678
rect 2389 638 2401 672
rect 2501 638 2513 672
rect 2389 632 2513 638
rect 2647 672 2771 678
rect 2647 638 2659 672
rect 2759 638 2771 672
rect 2647 632 2771 638
rect 2905 672 3029 678
rect 2905 638 2917 672
rect 3017 638 3029 672
rect 2905 632 3029 638
rect 3163 672 3287 678
rect 3163 638 3175 672
rect 3275 638 3287 672
rect 3163 632 3287 638
rect -3377 588 -3331 600
rect -3377 -588 -3371 588
rect -3337 -588 -3331 588
rect -3377 -600 -3331 -588
rect -3119 588 -3073 600
rect -3119 -588 -3113 588
rect -3079 -588 -3073 588
rect -3119 -600 -3073 -588
rect -2861 588 -2815 600
rect -2861 -588 -2855 588
rect -2821 -588 -2815 588
rect -2861 -600 -2815 -588
rect -2603 588 -2557 600
rect -2603 -588 -2597 588
rect -2563 -588 -2557 588
rect -2603 -600 -2557 -588
rect -2345 588 -2299 600
rect -2345 -588 -2339 588
rect -2305 -588 -2299 588
rect -2345 -600 -2299 -588
rect -2087 588 -2041 600
rect -2087 -588 -2081 588
rect -2047 -588 -2041 588
rect -2087 -600 -2041 -588
rect -1829 588 -1783 600
rect -1829 -588 -1823 588
rect -1789 -588 -1783 588
rect -1829 -600 -1783 -588
rect -1571 588 -1525 600
rect -1571 -588 -1565 588
rect -1531 -588 -1525 588
rect -1571 -600 -1525 -588
rect -1313 588 -1267 600
rect -1313 -588 -1307 588
rect -1273 -588 -1267 588
rect -1313 -600 -1267 -588
rect -1055 588 -1009 600
rect -1055 -588 -1049 588
rect -1015 -588 -1009 588
rect -1055 -600 -1009 -588
rect -797 588 -751 600
rect -797 -588 -791 588
rect -757 -588 -751 588
rect -797 -600 -751 -588
rect -539 588 -493 600
rect -539 -588 -533 588
rect -499 -588 -493 588
rect -539 -600 -493 -588
rect -281 588 -235 600
rect -281 -588 -275 588
rect -241 -588 -235 588
rect -281 -600 -235 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 235 588 281 600
rect 235 -588 241 588
rect 275 -588 281 588
rect 235 -600 281 -588
rect 493 588 539 600
rect 493 -588 499 588
rect 533 -588 539 588
rect 493 -600 539 -588
rect 751 588 797 600
rect 751 -588 757 588
rect 791 -588 797 588
rect 751 -600 797 -588
rect 1009 588 1055 600
rect 1009 -588 1015 588
rect 1049 -588 1055 588
rect 1009 -600 1055 -588
rect 1267 588 1313 600
rect 1267 -588 1273 588
rect 1307 -588 1313 588
rect 1267 -600 1313 -588
rect 1525 588 1571 600
rect 1525 -588 1531 588
rect 1565 -588 1571 588
rect 1525 -600 1571 -588
rect 1783 588 1829 600
rect 1783 -588 1789 588
rect 1823 -588 1829 588
rect 1783 -600 1829 -588
rect 2041 588 2087 600
rect 2041 -588 2047 588
rect 2081 -588 2087 588
rect 2041 -600 2087 -588
rect 2299 588 2345 600
rect 2299 -588 2305 588
rect 2339 -588 2345 588
rect 2299 -600 2345 -588
rect 2557 588 2603 600
rect 2557 -588 2563 588
rect 2597 -588 2603 588
rect 2557 -600 2603 -588
rect 2815 588 2861 600
rect 2815 -588 2821 588
rect 2855 -588 2861 588
rect 2815 -600 2861 -588
rect 3073 588 3119 600
rect 3073 -588 3079 588
rect 3113 -588 3119 588
rect 3073 -600 3119 -588
rect 3331 588 3377 600
rect 3331 -588 3337 588
rect 3371 -588 3377 588
rect 3331 -600 3377 -588
rect -3287 -638 -3163 -632
rect -3287 -672 -3275 -638
rect -3175 -672 -3163 -638
rect -3287 -678 -3163 -672
rect -3029 -638 -2905 -632
rect -3029 -672 -3017 -638
rect -2917 -672 -2905 -638
rect -3029 -678 -2905 -672
rect -2771 -638 -2647 -632
rect -2771 -672 -2759 -638
rect -2659 -672 -2647 -638
rect -2771 -678 -2647 -672
rect -2513 -638 -2389 -632
rect -2513 -672 -2501 -638
rect -2401 -672 -2389 -638
rect -2513 -678 -2389 -672
rect -2255 -638 -2131 -632
rect -2255 -672 -2243 -638
rect -2143 -672 -2131 -638
rect -2255 -678 -2131 -672
rect -1997 -638 -1873 -632
rect -1997 -672 -1985 -638
rect -1885 -672 -1873 -638
rect -1997 -678 -1873 -672
rect -1739 -638 -1615 -632
rect -1739 -672 -1727 -638
rect -1627 -672 -1615 -638
rect -1739 -678 -1615 -672
rect -1481 -638 -1357 -632
rect -1481 -672 -1469 -638
rect -1369 -672 -1357 -638
rect -1481 -678 -1357 -672
rect -1223 -638 -1099 -632
rect -1223 -672 -1211 -638
rect -1111 -672 -1099 -638
rect -1223 -678 -1099 -672
rect -965 -638 -841 -632
rect -965 -672 -953 -638
rect -853 -672 -841 -638
rect -965 -678 -841 -672
rect -707 -638 -583 -632
rect -707 -672 -695 -638
rect -595 -672 -583 -638
rect -707 -678 -583 -672
rect -449 -638 -325 -632
rect -449 -672 -437 -638
rect -337 -672 -325 -638
rect -449 -678 -325 -672
rect -191 -638 -67 -632
rect -191 -672 -179 -638
rect -79 -672 -67 -638
rect -191 -678 -67 -672
rect 67 -638 191 -632
rect 67 -672 79 -638
rect 179 -672 191 -638
rect 67 -678 191 -672
rect 325 -638 449 -632
rect 325 -672 337 -638
rect 437 -672 449 -638
rect 325 -678 449 -672
rect 583 -638 707 -632
rect 583 -672 595 -638
rect 695 -672 707 -638
rect 583 -678 707 -672
rect 841 -638 965 -632
rect 841 -672 853 -638
rect 953 -672 965 -638
rect 841 -678 965 -672
rect 1099 -638 1223 -632
rect 1099 -672 1111 -638
rect 1211 -672 1223 -638
rect 1099 -678 1223 -672
rect 1357 -638 1481 -632
rect 1357 -672 1369 -638
rect 1469 -672 1481 -638
rect 1357 -678 1481 -672
rect 1615 -638 1739 -632
rect 1615 -672 1627 -638
rect 1727 -672 1739 -638
rect 1615 -678 1739 -672
rect 1873 -638 1997 -632
rect 1873 -672 1885 -638
rect 1985 -672 1997 -638
rect 1873 -678 1997 -672
rect 2131 -638 2255 -632
rect 2131 -672 2143 -638
rect 2243 -672 2255 -638
rect 2131 -678 2255 -672
rect 2389 -638 2513 -632
rect 2389 -672 2401 -638
rect 2501 -672 2513 -638
rect 2389 -678 2513 -672
rect 2647 -638 2771 -632
rect 2647 -672 2659 -638
rect 2759 -672 2771 -638
rect 2647 -678 2771 -672
rect 2905 -638 3029 -632
rect 2905 -672 2917 -638
rect 3017 -672 3029 -638
rect 2905 -678 3029 -672
rect 3163 -638 3287 -632
rect 3163 -672 3175 -638
rect 3275 -672 3287 -638
rect 3163 -678 3287 -672
<< properties >>
string FIXED_BBOX -3488 -793 3488 793
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6 l 1 m 1 nf 26 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713232286
<< pwell >>
rect -3553 -967 3553 967
<< mvnmos >>
rect -3325 109 -3125 709
rect -3067 109 -2867 709
rect -2809 109 -2609 709
rect -2551 109 -2351 709
rect -2293 109 -2093 709
rect -2035 109 -1835 709
rect -1777 109 -1577 709
rect -1519 109 -1319 709
rect -1261 109 -1061 709
rect -1003 109 -803 709
rect -745 109 -545 709
rect -487 109 -287 709
rect -229 109 -29 709
rect 29 109 229 709
rect 287 109 487 709
rect 545 109 745 709
rect 803 109 1003 709
rect 1061 109 1261 709
rect 1319 109 1519 709
rect 1577 109 1777 709
rect 1835 109 2035 709
rect 2093 109 2293 709
rect 2351 109 2551 709
rect 2609 109 2809 709
rect 2867 109 3067 709
rect 3125 109 3325 709
rect -3325 -709 -3125 -109
rect -3067 -709 -2867 -109
rect -2809 -709 -2609 -109
rect -2551 -709 -2351 -109
rect -2293 -709 -2093 -109
rect -2035 -709 -1835 -109
rect -1777 -709 -1577 -109
rect -1519 -709 -1319 -109
rect -1261 -709 -1061 -109
rect -1003 -709 -803 -109
rect -745 -709 -545 -109
rect -487 -709 -287 -109
rect -229 -709 -29 -109
rect 29 -709 229 -109
rect 287 -709 487 -109
rect 545 -709 745 -109
rect 803 -709 1003 -109
rect 1061 -709 1261 -109
rect 1319 -709 1519 -109
rect 1577 -709 1777 -109
rect 1835 -709 2035 -109
rect 2093 -709 2293 -109
rect 2351 -709 2551 -109
rect 2609 -709 2809 -109
rect 2867 -709 3067 -109
rect 3125 -709 3325 -109
<< mvndiff >>
rect -3383 697 -3325 709
rect -3383 121 -3371 697
rect -3337 121 -3325 697
rect -3383 109 -3325 121
rect -3125 697 -3067 709
rect -3125 121 -3113 697
rect -3079 121 -3067 697
rect -3125 109 -3067 121
rect -2867 697 -2809 709
rect -2867 121 -2855 697
rect -2821 121 -2809 697
rect -2867 109 -2809 121
rect -2609 697 -2551 709
rect -2609 121 -2597 697
rect -2563 121 -2551 697
rect -2609 109 -2551 121
rect -2351 697 -2293 709
rect -2351 121 -2339 697
rect -2305 121 -2293 697
rect -2351 109 -2293 121
rect -2093 697 -2035 709
rect -2093 121 -2081 697
rect -2047 121 -2035 697
rect -2093 109 -2035 121
rect -1835 697 -1777 709
rect -1835 121 -1823 697
rect -1789 121 -1777 697
rect -1835 109 -1777 121
rect -1577 697 -1519 709
rect -1577 121 -1565 697
rect -1531 121 -1519 697
rect -1577 109 -1519 121
rect -1319 697 -1261 709
rect -1319 121 -1307 697
rect -1273 121 -1261 697
rect -1319 109 -1261 121
rect -1061 697 -1003 709
rect -1061 121 -1049 697
rect -1015 121 -1003 697
rect -1061 109 -1003 121
rect -803 697 -745 709
rect -803 121 -791 697
rect -757 121 -745 697
rect -803 109 -745 121
rect -545 697 -487 709
rect -545 121 -533 697
rect -499 121 -487 697
rect -545 109 -487 121
rect -287 697 -229 709
rect -287 121 -275 697
rect -241 121 -229 697
rect -287 109 -229 121
rect -29 697 29 709
rect -29 121 -17 697
rect 17 121 29 697
rect -29 109 29 121
rect 229 697 287 709
rect 229 121 241 697
rect 275 121 287 697
rect 229 109 287 121
rect 487 697 545 709
rect 487 121 499 697
rect 533 121 545 697
rect 487 109 545 121
rect 745 697 803 709
rect 745 121 757 697
rect 791 121 803 697
rect 745 109 803 121
rect 1003 697 1061 709
rect 1003 121 1015 697
rect 1049 121 1061 697
rect 1003 109 1061 121
rect 1261 697 1319 709
rect 1261 121 1273 697
rect 1307 121 1319 697
rect 1261 109 1319 121
rect 1519 697 1577 709
rect 1519 121 1531 697
rect 1565 121 1577 697
rect 1519 109 1577 121
rect 1777 697 1835 709
rect 1777 121 1789 697
rect 1823 121 1835 697
rect 1777 109 1835 121
rect 2035 697 2093 709
rect 2035 121 2047 697
rect 2081 121 2093 697
rect 2035 109 2093 121
rect 2293 697 2351 709
rect 2293 121 2305 697
rect 2339 121 2351 697
rect 2293 109 2351 121
rect 2551 697 2609 709
rect 2551 121 2563 697
rect 2597 121 2609 697
rect 2551 109 2609 121
rect 2809 697 2867 709
rect 2809 121 2821 697
rect 2855 121 2867 697
rect 2809 109 2867 121
rect 3067 697 3125 709
rect 3067 121 3079 697
rect 3113 121 3125 697
rect 3067 109 3125 121
rect 3325 697 3383 709
rect 3325 121 3337 697
rect 3371 121 3383 697
rect 3325 109 3383 121
rect -3383 -121 -3325 -109
rect -3383 -697 -3371 -121
rect -3337 -697 -3325 -121
rect -3383 -709 -3325 -697
rect -3125 -121 -3067 -109
rect -3125 -697 -3113 -121
rect -3079 -697 -3067 -121
rect -3125 -709 -3067 -697
rect -2867 -121 -2809 -109
rect -2867 -697 -2855 -121
rect -2821 -697 -2809 -121
rect -2867 -709 -2809 -697
rect -2609 -121 -2551 -109
rect -2609 -697 -2597 -121
rect -2563 -697 -2551 -121
rect -2609 -709 -2551 -697
rect -2351 -121 -2293 -109
rect -2351 -697 -2339 -121
rect -2305 -697 -2293 -121
rect -2351 -709 -2293 -697
rect -2093 -121 -2035 -109
rect -2093 -697 -2081 -121
rect -2047 -697 -2035 -121
rect -2093 -709 -2035 -697
rect -1835 -121 -1777 -109
rect -1835 -697 -1823 -121
rect -1789 -697 -1777 -121
rect -1835 -709 -1777 -697
rect -1577 -121 -1519 -109
rect -1577 -697 -1565 -121
rect -1531 -697 -1519 -121
rect -1577 -709 -1519 -697
rect -1319 -121 -1261 -109
rect -1319 -697 -1307 -121
rect -1273 -697 -1261 -121
rect -1319 -709 -1261 -697
rect -1061 -121 -1003 -109
rect -1061 -697 -1049 -121
rect -1015 -697 -1003 -121
rect -1061 -709 -1003 -697
rect -803 -121 -745 -109
rect -803 -697 -791 -121
rect -757 -697 -745 -121
rect -803 -709 -745 -697
rect -545 -121 -487 -109
rect -545 -697 -533 -121
rect -499 -697 -487 -121
rect -545 -709 -487 -697
rect -287 -121 -229 -109
rect -287 -697 -275 -121
rect -241 -697 -229 -121
rect -287 -709 -229 -697
rect -29 -121 29 -109
rect -29 -697 -17 -121
rect 17 -697 29 -121
rect -29 -709 29 -697
rect 229 -121 287 -109
rect 229 -697 241 -121
rect 275 -697 287 -121
rect 229 -709 287 -697
rect 487 -121 545 -109
rect 487 -697 499 -121
rect 533 -697 545 -121
rect 487 -709 545 -697
rect 745 -121 803 -109
rect 745 -697 757 -121
rect 791 -697 803 -121
rect 745 -709 803 -697
rect 1003 -121 1061 -109
rect 1003 -697 1015 -121
rect 1049 -697 1061 -121
rect 1003 -709 1061 -697
rect 1261 -121 1319 -109
rect 1261 -697 1273 -121
rect 1307 -697 1319 -121
rect 1261 -709 1319 -697
rect 1519 -121 1577 -109
rect 1519 -697 1531 -121
rect 1565 -697 1577 -121
rect 1519 -709 1577 -697
rect 1777 -121 1835 -109
rect 1777 -697 1789 -121
rect 1823 -697 1835 -121
rect 1777 -709 1835 -697
rect 2035 -121 2093 -109
rect 2035 -697 2047 -121
rect 2081 -697 2093 -121
rect 2035 -709 2093 -697
rect 2293 -121 2351 -109
rect 2293 -697 2305 -121
rect 2339 -697 2351 -121
rect 2293 -709 2351 -697
rect 2551 -121 2609 -109
rect 2551 -697 2563 -121
rect 2597 -697 2609 -121
rect 2551 -709 2609 -697
rect 2809 -121 2867 -109
rect 2809 -697 2821 -121
rect 2855 -697 2867 -121
rect 2809 -709 2867 -697
rect 3067 -121 3125 -109
rect 3067 -697 3079 -121
rect 3113 -697 3125 -121
rect 3067 -709 3125 -697
rect 3325 -121 3383 -109
rect 3325 -697 3337 -121
rect 3371 -697 3383 -121
rect 3325 -709 3383 -697
<< mvndiffc >>
rect -3371 121 -3337 697
rect -3113 121 -3079 697
rect -2855 121 -2821 697
rect -2597 121 -2563 697
rect -2339 121 -2305 697
rect -2081 121 -2047 697
rect -1823 121 -1789 697
rect -1565 121 -1531 697
rect -1307 121 -1273 697
rect -1049 121 -1015 697
rect -791 121 -757 697
rect -533 121 -499 697
rect -275 121 -241 697
rect -17 121 17 697
rect 241 121 275 697
rect 499 121 533 697
rect 757 121 791 697
rect 1015 121 1049 697
rect 1273 121 1307 697
rect 1531 121 1565 697
rect 1789 121 1823 697
rect 2047 121 2081 697
rect 2305 121 2339 697
rect 2563 121 2597 697
rect 2821 121 2855 697
rect 3079 121 3113 697
rect 3337 121 3371 697
rect -3371 -697 -3337 -121
rect -3113 -697 -3079 -121
rect -2855 -697 -2821 -121
rect -2597 -697 -2563 -121
rect -2339 -697 -2305 -121
rect -2081 -697 -2047 -121
rect -1823 -697 -1789 -121
rect -1565 -697 -1531 -121
rect -1307 -697 -1273 -121
rect -1049 -697 -1015 -121
rect -791 -697 -757 -121
rect -533 -697 -499 -121
rect -275 -697 -241 -121
rect -17 -697 17 -121
rect 241 -697 275 -121
rect 499 -697 533 -121
rect 757 -697 791 -121
rect 1015 -697 1049 -121
rect 1273 -697 1307 -121
rect 1531 -697 1565 -121
rect 1789 -697 1823 -121
rect 2047 -697 2081 -121
rect 2305 -697 2339 -121
rect 2563 -697 2597 -121
rect 2821 -697 2855 -121
rect 3079 -697 3113 -121
rect 3337 -697 3371 -121
<< mvpsubdiff >>
rect -3517 919 3517 931
rect -3517 885 -3409 919
rect 3409 885 3517 919
rect -3517 873 3517 885
rect -3517 823 -3459 873
rect -3517 -823 -3505 823
rect -3471 -823 -3459 823
rect 3459 823 3517 873
rect -3517 -873 -3459 -823
rect 3459 -823 3471 823
rect 3505 -823 3517 823
rect 3459 -873 3517 -823
rect -3517 -885 3517 -873
rect -3517 -919 -3409 -885
rect 3409 -919 3517 -885
rect -3517 -931 3517 -919
<< mvpsubdiffcont >>
rect -3409 885 3409 919
rect -3505 -823 -3471 823
rect 3471 -823 3505 823
rect -3409 -919 3409 -885
<< poly >>
rect -3325 781 -3125 797
rect -3325 747 -3309 781
rect -3141 747 -3125 781
rect -3325 709 -3125 747
rect -3067 781 -2867 797
rect -3067 747 -3051 781
rect -2883 747 -2867 781
rect -3067 709 -2867 747
rect -2809 781 -2609 797
rect -2809 747 -2793 781
rect -2625 747 -2609 781
rect -2809 709 -2609 747
rect -2551 781 -2351 797
rect -2551 747 -2535 781
rect -2367 747 -2351 781
rect -2551 709 -2351 747
rect -2293 781 -2093 797
rect -2293 747 -2277 781
rect -2109 747 -2093 781
rect -2293 709 -2093 747
rect -2035 781 -1835 797
rect -2035 747 -2019 781
rect -1851 747 -1835 781
rect -2035 709 -1835 747
rect -1777 781 -1577 797
rect -1777 747 -1761 781
rect -1593 747 -1577 781
rect -1777 709 -1577 747
rect -1519 781 -1319 797
rect -1519 747 -1503 781
rect -1335 747 -1319 781
rect -1519 709 -1319 747
rect -1261 781 -1061 797
rect -1261 747 -1245 781
rect -1077 747 -1061 781
rect -1261 709 -1061 747
rect -1003 781 -803 797
rect -1003 747 -987 781
rect -819 747 -803 781
rect -1003 709 -803 747
rect -745 781 -545 797
rect -745 747 -729 781
rect -561 747 -545 781
rect -745 709 -545 747
rect -487 781 -287 797
rect -487 747 -471 781
rect -303 747 -287 781
rect -487 709 -287 747
rect -229 781 -29 797
rect -229 747 -213 781
rect -45 747 -29 781
rect -229 709 -29 747
rect 29 781 229 797
rect 29 747 45 781
rect 213 747 229 781
rect 29 709 229 747
rect 287 781 487 797
rect 287 747 303 781
rect 471 747 487 781
rect 287 709 487 747
rect 545 781 745 797
rect 545 747 561 781
rect 729 747 745 781
rect 545 709 745 747
rect 803 781 1003 797
rect 803 747 819 781
rect 987 747 1003 781
rect 803 709 1003 747
rect 1061 781 1261 797
rect 1061 747 1077 781
rect 1245 747 1261 781
rect 1061 709 1261 747
rect 1319 781 1519 797
rect 1319 747 1335 781
rect 1503 747 1519 781
rect 1319 709 1519 747
rect 1577 781 1777 797
rect 1577 747 1593 781
rect 1761 747 1777 781
rect 1577 709 1777 747
rect 1835 781 2035 797
rect 1835 747 1851 781
rect 2019 747 2035 781
rect 1835 709 2035 747
rect 2093 781 2293 797
rect 2093 747 2109 781
rect 2277 747 2293 781
rect 2093 709 2293 747
rect 2351 781 2551 797
rect 2351 747 2367 781
rect 2535 747 2551 781
rect 2351 709 2551 747
rect 2609 781 2809 797
rect 2609 747 2625 781
rect 2793 747 2809 781
rect 2609 709 2809 747
rect 2867 781 3067 797
rect 2867 747 2883 781
rect 3051 747 3067 781
rect 2867 709 3067 747
rect 3125 781 3325 797
rect 3125 747 3141 781
rect 3309 747 3325 781
rect 3125 709 3325 747
rect -3325 71 -3125 109
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3325 21 -3125 37
rect -3067 71 -2867 109
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -3067 21 -2867 37
rect -2809 71 -2609 109
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2809 21 -2609 37
rect -2551 71 -2351 109
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2551 21 -2351 37
rect -2293 71 -2093 109
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2293 21 -2093 37
rect -2035 71 -1835 109
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 109
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 109
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 109
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 109
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 109
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 109
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 109
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 109
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 109
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 109
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 109
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 109
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 109
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 109
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 109
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect 2093 71 2293 109
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2093 21 2293 37
rect 2351 71 2551 109
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2351 21 2551 37
rect 2609 71 2809 109
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2609 21 2809 37
rect 2867 71 3067 109
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 2867 21 3067 37
rect 3125 71 3325 109
rect 3125 37 3141 71
rect 3309 37 3325 71
rect 3125 21 3325 37
rect -3325 -37 -3125 -21
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3325 -109 -3125 -71
rect -3067 -37 -2867 -21
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -3067 -109 -2867 -71
rect -2809 -37 -2609 -21
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2809 -109 -2609 -71
rect -2551 -37 -2351 -21
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2551 -109 -2351 -71
rect -2293 -37 -2093 -21
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2293 -109 -2093 -71
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -109 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -109 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -109 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -109 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -109 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -109 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -109 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -109 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -109 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -109 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -109 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -109 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -109 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -109 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -109 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -109 2035 -71
rect 2093 -37 2293 -21
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2093 -109 2293 -71
rect 2351 -37 2551 -21
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2351 -109 2551 -71
rect 2609 -37 2809 -21
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2609 -109 2809 -71
rect 2867 -37 3067 -21
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 2867 -109 3067 -71
rect 3125 -37 3325 -21
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect 3125 -109 3325 -71
rect -3325 -747 -3125 -709
rect -3325 -781 -3309 -747
rect -3141 -781 -3125 -747
rect -3325 -797 -3125 -781
rect -3067 -747 -2867 -709
rect -3067 -781 -3051 -747
rect -2883 -781 -2867 -747
rect -3067 -797 -2867 -781
rect -2809 -747 -2609 -709
rect -2809 -781 -2793 -747
rect -2625 -781 -2609 -747
rect -2809 -797 -2609 -781
rect -2551 -747 -2351 -709
rect -2551 -781 -2535 -747
rect -2367 -781 -2351 -747
rect -2551 -797 -2351 -781
rect -2293 -747 -2093 -709
rect -2293 -781 -2277 -747
rect -2109 -781 -2093 -747
rect -2293 -797 -2093 -781
rect -2035 -747 -1835 -709
rect -2035 -781 -2019 -747
rect -1851 -781 -1835 -747
rect -2035 -797 -1835 -781
rect -1777 -747 -1577 -709
rect -1777 -781 -1761 -747
rect -1593 -781 -1577 -747
rect -1777 -797 -1577 -781
rect -1519 -747 -1319 -709
rect -1519 -781 -1503 -747
rect -1335 -781 -1319 -747
rect -1519 -797 -1319 -781
rect -1261 -747 -1061 -709
rect -1261 -781 -1245 -747
rect -1077 -781 -1061 -747
rect -1261 -797 -1061 -781
rect -1003 -747 -803 -709
rect -1003 -781 -987 -747
rect -819 -781 -803 -747
rect -1003 -797 -803 -781
rect -745 -747 -545 -709
rect -745 -781 -729 -747
rect -561 -781 -545 -747
rect -745 -797 -545 -781
rect -487 -747 -287 -709
rect -487 -781 -471 -747
rect -303 -781 -287 -747
rect -487 -797 -287 -781
rect -229 -747 -29 -709
rect -229 -781 -213 -747
rect -45 -781 -29 -747
rect -229 -797 -29 -781
rect 29 -747 229 -709
rect 29 -781 45 -747
rect 213 -781 229 -747
rect 29 -797 229 -781
rect 287 -747 487 -709
rect 287 -781 303 -747
rect 471 -781 487 -747
rect 287 -797 487 -781
rect 545 -747 745 -709
rect 545 -781 561 -747
rect 729 -781 745 -747
rect 545 -797 745 -781
rect 803 -747 1003 -709
rect 803 -781 819 -747
rect 987 -781 1003 -747
rect 803 -797 1003 -781
rect 1061 -747 1261 -709
rect 1061 -781 1077 -747
rect 1245 -781 1261 -747
rect 1061 -797 1261 -781
rect 1319 -747 1519 -709
rect 1319 -781 1335 -747
rect 1503 -781 1519 -747
rect 1319 -797 1519 -781
rect 1577 -747 1777 -709
rect 1577 -781 1593 -747
rect 1761 -781 1777 -747
rect 1577 -797 1777 -781
rect 1835 -747 2035 -709
rect 1835 -781 1851 -747
rect 2019 -781 2035 -747
rect 1835 -797 2035 -781
rect 2093 -747 2293 -709
rect 2093 -781 2109 -747
rect 2277 -781 2293 -747
rect 2093 -797 2293 -781
rect 2351 -747 2551 -709
rect 2351 -781 2367 -747
rect 2535 -781 2551 -747
rect 2351 -797 2551 -781
rect 2609 -747 2809 -709
rect 2609 -781 2625 -747
rect 2793 -781 2809 -747
rect 2609 -797 2809 -781
rect 2867 -747 3067 -709
rect 2867 -781 2883 -747
rect 3051 -781 3067 -747
rect 2867 -797 3067 -781
rect 3125 -747 3325 -709
rect 3125 -781 3141 -747
rect 3309 -781 3325 -747
rect 3125 -797 3325 -781
<< polycont >>
rect -3309 747 -3141 781
rect -3051 747 -2883 781
rect -2793 747 -2625 781
rect -2535 747 -2367 781
rect -2277 747 -2109 781
rect -2019 747 -1851 781
rect -1761 747 -1593 781
rect -1503 747 -1335 781
rect -1245 747 -1077 781
rect -987 747 -819 781
rect -729 747 -561 781
rect -471 747 -303 781
rect -213 747 -45 781
rect 45 747 213 781
rect 303 747 471 781
rect 561 747 729 781
rect 819 747 987 781
rect 1077 747 1245 781
rect 1335 747 1503 781
rect 1593 747 1761 781
rect 1851 747 2019 781
rect 2109 747 2277 781
rect 2367 747 2535 781
rect 2625 747 2793 781
rect 2883 747 3051 781
rect 3141 747 3309 781
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect -3309 -781 -3141 -747
rect -3051 -781 -2883 -747
rect -2793 -781 -2625 -747
rect -2535 -781 -2367 -747
rect -2277 -781 -2109 -747
rect -2019 -781 -1851 -747
rect -1761 -781 -1593 -747
rect -1503 -781 -1335 -747
rect -1245 -781 -1077 -747
rect -987 -781 -819 -747
rect -729 -781 -561 -747
rect -471 -781 -303 -747
rect -213 -781 -45 -747
rect 45 -781 213 -747
rect 303 -781 471 -747
rect 561 -781 729 -747
rect 819 -781 987 -747
rect 1077 -781 1245 -747
rect 1335 -781 1503 -747
rect 1593 -781 1761 -747
rect 1851 -781 2019 -747
rect 2109 -781 2277 -747
rect 2367 -781 2535 -747
rect 2625 -781 2793 -747
rect 2883 -781 3051 -747
rect 3141 -781 3309 -747
<< locali >>
rect -3505 885 -3409 919
rect 3409 885 3505 919
rect -3505 823 -3471 885
rect 3471 823 3505 885
rect -3325 747 -3309 781
rect -3141 747 -3125 781
rect -3067 747 -3051 781
rect -2883 747 -2867 781
rect -2809 747 -2793 781
rect -2625 747 -2609 781
rect -2551 747 -2535 781
rect -2367 747 -2351 781
rect -2293 747 -2277 781
rect -2109 747 -2093 781
rect -2035 747 -2019 781
rect -1851 747 -1835 781
rect -1777 747 -1761 781
rect -1593 747 -1577 781
rect -1519 747 -1503 781
rect -1335 747 -1319 781
rect -1261 747 -1245 781
rect -1077 747 -1061 781
rect -1003 747 -987 781
rect -819 747 -803 781
rect -745 747 -729 781
rect -561 747 -545 781
rect -487 747 -471 781
rect -303 747 -287 781
rect -229 747 -213 781
rect -45 747 -29 781
rect 29 747 45 781
rect 213 747 229 781
rect 287 747 303 781
rect 471 747 487 781
rect 545 747 561 781
rect 729 747 745 781
rect 803 747 819 781
rect 987 747 1003 781
rect 1061 747 1077 781
rect 1245 747 1261 781
rect 1319 747 1335 781
rect 1503 747 1519 781
rect 1577 747 1593 781
rect 1761 747 1777 781
rect 1835 747 1851 781
rect 2019 747 2035 781
rect 2093 747 2109 781
rect 2277 747 2293 781
rect 2351 747 2367 781
rect 2535 747 2551 781
rect 2609 747 2625 781
rect 2793 747 2809 781
rect 2867 747 2883 781
rect 3051 747 3067 781
rect 3125 747 3141 781
rect 3309 747 3325 781
rect -3371 697 -3337 713
rect -3371 105 -3337 121
rect -3113 697 -3079 713
rect -3113 105 -3079 121
rect -2855 697 -2821 713
rect -2855 105 -2821 121
rect -2597 697 -2563 713
rect -2597 105 -2563 121
rect -2339 697 -2305 713
rect -2339 105 -2305 121
rect -2081 697 -2047 713
rect -2081 105 -2047 121
rect -1823 697 -1789 713
rect -1823 105 -1789 121
rect -1565 697 -1531 713
rect -1565 105 -1531 121
rect -1307 697 -1273 713
rect -1307 105 -1273 121
rect -1049 697 -1015 713
rect -1049 105 -1015 121
rect -791 697 -757 713
rect -791 105 -757 121
rect -533 697 -499 713
rect -533 105 -499 121
rect -275 697 -241 713
rect -275 105 -241 121
rect -17 697 17 713
rect -17 105 17 121
rect 241 697 275 713
rect 241 105 275 121
rect 499 697 533 713
rect 499 105 533 121
rect 757 697 791 713
rect 757 105 791 121
rect 1015 697 1049 713
rect 1015 105 1049 121
rect 1273 697 1307 713
rect 1273 105 1307 121
rect 1531 697 1565 713
rect 1531 105 1565 121
rect 1789 697 1823 713
rect 1789 105 1823 121
rect 2047 697 2081 713
rect 2047 105 2081 121
rect 2305 697 2339 713
rect 2305 105 2339 121
rect 2563 697 2597 713
rect 2563 105 2597 121
rect 2821 697 2855 713
rect 2821 105 2855 121
rect 3079 697 3113 713
rect 3079 105 3113 121
rect 3337 697 3371 713
rect 3337 105 3371 121
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 3125 37 3141 71
rect 3309 37 3325 71
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect -3371 -121 -3337 -105
rect -3371 -713 -3337 -697
rect -3113 -121 -3079 -105
rect -3113 -713 -3079 -697
rect -2855 -121 -2821 -105
rect -2855 -713 -2821 -697
rect -2597 -121 -2563 -105
rect -2597 -713 -2563 -697
rect -2339 -121 -2305 -105
rect -2339 -713 -2305 -697
rect -2081 -121 -2047 -105
rect -2081 -713 -2047 -697
rect -1823 -121 -1789 -105
rect -1823 -713 -1789 -697
rect -1565 -121 -1531 -105
rect -1565 -713 -1531 -697
rect -1307 -121 -1273 -105
rect -1307 -713 -1273 -697
rect -1049 -121 -1015 -105
rect -1049 -713 -1015 -697
rect -791 -121 -757 -105
rect -791 -713 -757 -697
rect -533 -121 -499 -105
rect -533 -713 -499 -697
rect -275 -121 -241 -105
rect -275 -713 -241 -697
rect -17 -121 17 -105
rect -17 -713 17 -697
rect 241 -121 275 -105
rect 241 -713 275 -697
rect 499 -121 533 -105
rect 499 -713 533 -697
rect 757 -121 791 -105
rect 757 -713 791 -697
rect 1015 -121 1049 -105
rect 1015 -713 1049 -697
rect 1273 -121 1307 -105
rect 1273 -713 1307 -697
rect 1531 -121 1565 -105
rect 1531 -713 1565 -697
rect 1789 -121 1823 -105
rect 1789 -713 1823 -697
rect 2047 -121 2081 -105
rect 2047 -713 2081 -697
rect 2305 -121 2339 -105
rect 2305 -713 2339 -697
rect 2563 -121 2597 -105
rect 2563 -713 2597 -697
rect 2821 -121 2855 -105
rect 2821 -713 2855 -697
rect 3079 -121 3113 -105
rect 3079 -713 3113 -697
rect 3337 -121 3371 -105
rect 3337 -713 3371 -697
rect -3325 -781 -3309 -747
rect -3141 -781 -3125 -747
rect -3067 -781 -3051 -747
rect -2883 -781 -2867 -747
rect -2809 -781 -2793 -747
rect -2625 -781 -2609 -747
rect -2551 -781 -2535 -747
rect -2367 -781 -2351 -747
rect -2293 -781 -2277 -747
rect -2109 -781 -2093 -747
rect -2035 -781 -2019 -747
rect -1851 -781 -1835 -747
rect -1777 -781 -1761 -747
rect -1593 -781 -1577 -747
rect -1519 -781 -1503 -747
rect -1335 -781 -1319 -747
rect -1261 -781 -1245 -747
rect -1077 -781 -1061 -747
rect -1003 -781 -987 -747
rect -819 -781 -803 -747
rect -745 -781 -729 -747
rect -561 -781 -545 -747
rect -487 -781 -471 -747
rect -303 -781 -287 -747
rect -229 -781 -213 -747
rect -45 -781 -29 -747
rect 29 -781 45 -747
rect 213 -781 229 -747
rect 287 -781 303 -747
rect 471 -781 487 -747
rect 545 -781 561 -747
rect 729 -781 745 -747
rect 803 -781 819 -747
rect 987 -781 1003 -747
rect 1061 -781 1077 -747
rect 1245 -781 1261 -747
rect 1319 -781 1335 -747
rect 1503 -781 1519 -747
rect 1577 -781 1593 -747
rect 1761 -781 1777 -747
rect 1835 -781 1851 -747
rect 2019 -781 2035 -747
rect 2093 -781 2109 -747
rect 2277 -781 2293 -747
rect 2351 -781 2367 -747
rect 2535 -781 2551 -747
rect 2609 -781 2625 -747
rect 2793 -781 2809 -747
rect 2867 -781 2883 -747
rect 3051 -781 3067 -747
rect 3125 -781 3141 -747
rect 3309 -781 3325 -747
rect -3505 -885 -3471 -823
rect 3471 -885 3505 -823
rect -3505 -919 -3409 -885
rect 3409 -919 3505 -885
<< viali >>
rect -3309 747 -3141 781
rect -3051 747 -2883 781
rect -2793 747 -2625 781
rect -2535 747 -2367 781
rect -2277 747 -2109 781
rect -2019 747 -1851 781
rect -1761 747 -1593 781
rect -1503 747 -1335 781
rect -1245 747 -1077 781
rect -987 747 -819 781
rect -729 747 -561 781
rect -471 747 -303 781
rect -213 747 -45 781
rect 45 747 213 781
rect 303 747 471 781
rect 561 747 729 781
rect 819 747 987 781
rect 1077 747 1245 781
rect 1335 747 1503 781
rect 1593 747 1761 781
rect 1851 747 2019 781
rect 2109 747 2277 781
rect 2367 747 2535 781
rect 2625 747 2793 781
rect 2883 747 3051 781
rect 3141 747 3309 781
rect -3371 121 -3337 697
rect -3113 121 -3079 697
rect -2855 121 -2821 697
rect -2597 121 -2563 697
rect -2339 121 -2305 697
rect -2081 121 -2047 697
rect -1823 121 -1789 697
rect -1565 121 -1531 697
rect -1307 121 -1273 697
rect -1049 121 -1015 697
rect -791 121 -757 697
rect -533 121 -499 697
rect -275 121 -241 697
rect -17 121 17 697
rect 241 121 275 697
rect 499 121 533 697
rect 757 121 791 697
rect 1015 121 1049 697
rect 1273 121 1307 697
rect 1531 121 1565 697
rect 1789 121 1823 697
rect 2047 121 2081 697
rect 2305 121 2339 697
rect 2563 121 2597 697
rect 2821 121 2855 697
rect 3079 121 3113 697
rect 3337 121 3371 697
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect -3371 -697 -3337 -121
rect -3113 -697 -3079 -121
rect -2855 -697 -2821 -121
rect -2597 -697 -2563 -121
rect -2339 -697 -2305 -121
rect -2081 -697 -2047 -121
rect -1823 -697 -1789 -121
rect -1565 -697 -1531 -121
rect -1307 -697 -1273 -121
rect -1049 -697 -1015 -121
rect -791 -697 -757 -121
rect -533 -697 -499 -121
rect -275 -697 -241 -121
rect -17 -697 17 -121
rect 241 -697 275 -121
rect 499 -697 533 -121
rect 757 -697 791 -121
rect 1015 -697 1049 -121
rect 1273 -697 1307 -121
rect 1531 -697 1565 -121
rect 1789 -697 1823 -121
rect 2047 -697 2081 -121
rect 2305 -697 2339 -121
rect 2563 -697 2597 -121
rect 2821 -697 2855 -121
rect 3079 -697 3113 -121
rect 3337 -697 3371 -121
rect -3309 -781 -3141 -747
rect -3051 -781 -2883 -747
rect -2793 -781 -2625 -747
rect -2535 -781 -2367 -747
rect -2277 -781 -2109 -747
rect -2019 -781 -1851 -747
rect -1761 -781 -1593 -747
rect -1503 -781 -1335 -747
rect -1245 -781 -1077 -747
rect -987 -781 -819 -747
rect -729 -781 -561 -747
rect -471 -781 -303 -747
rect -213 -781 -45 -747
rect 45 -781 213 -747
rect 303 -781 471 -747
rect 561 -781 729 -747
rect 819 -781 987 -747
rect 1077 -781 1245 -747
rect 1335 -781 1503 -747
rect 1593 -781 1761 -747
rect 1851 -781 2019 -747
rect 2109 -781 2277 -747
rect 2367 -781 2535 -747
rect 2625 -781 2793 -747
rect 2883 -781 3051 -747
rect 3141 -781 3309 -747
<< metal1 >>
rect -3321 781 -3129 787
rect -3321 747 -3309 781
rect -3141 747 -3129 781
rect -3321 741 -3129 747
rect -3063 781 -2871 787
rect -3063 747 -3051 781
rect -2883 747 -2871 781
rect -3063 741 -2871 747
rect -2805 781 -2613 787
rect -2805 747 -2793 781
rect -2625 747 -2613 781
rect -2805 741 -2613 747
rect -2547 781 -2355 787
rect -2547 747 -2535 781
rect -2367 747 -2355 781
rect -2547 741 -2355 747
rect -2289 781 -2097 787
rect -2289 747 -2277 781
rect -2109 747 -2097 781
rect -2289 741 -2097 747
rect -2031 781 -1839 787
rect -2031 747 -2019 781
rect -1851 747 -1839 781
rect -2031 741 -1839 747
rect -1773 781 -1581 787
rect -1773 747 -1761 781
rect -1593 747 -1581 781
rect -1773 741 -1581 747
rect -1515 781 -1323 787
rect -1515 747 -1503 781
rect -1335 747 -1323 781
rect -1515 741 -1323 747
rect -1257 781 -1065 787
rect -1257 747 -1245 781
rect -1077 747 -1065 781
rect -1257 741 -1065 747
rect -999 781 -807 787
rect -999 747 -987 781
rect -819 747 -807 781
rect -999 741 -807 747
rect -741 781 -549 787
rect -741 747 -729 781
rect -561 747 -549 781
rect -741 741 -549 747
rect -483 781 -291 787
rect -483 747 -471 781
rect -303 747 -291 781
rect -483 741 -291 747
rect -225 781 -33 787
rect -225 747 -213 781
rect -45 747 -33 781
rect -225 741 -33 747
rect 33 781 225 787
rect 33 747 45 781
rect 213 747 225 781
rect 33 741 225 747
rect 291 781 483 787
rect 291 747 303 781
rect 471 747 483 781
rect 291 741 483 747
rect 549 781 741 787
rect 549 747 561 781
rect 729 747 741 781
rect 549 741 741 747
rect 807 781 999 787
rect 807 747 819 781
rect 987 747 999 781
rect 807 741 999 747
rect 1065 781 1257 787
rect 1065 747 1077 781
rect 1245 747 1257 781
rect 1065 741 1257 747
rect 1323 781 1515 787
rect 1323 747 1335 781
rect 1503 747 1515 781
rect 1323 741 1515 747
rect 1581 781 1773 787
rect 1581 747 1593 781
rect 1761 747 1773 781
rect 1581 741 1773 747
rect 1839 781 2031 787
rect 1839 747 1851 781
rect 2019 747 2031 781
rect 1839 741 2031 747
rect 2097 781 2289 787
rect 2097 747 2109 781
rect 2277 747 2289 781
rect 2097 741 2289 747
rect 2355 781 2547 787
rect 2355 747 2367 781
rect 2535 747 2547 781
rect 2355 741 2547 747
rect 2613 781 2805 787
rect 2613 747 2625 781
rect 2793 747 2805 781
rect 2613 741 2805 747
rect 2871 781 3063 787
rect 2871 747 2883 781
rect 3051 747 3063 781
rect 2871 741 3063 747
rect 3129 781 3321 787
rect 3129 747 3141 781
rect 3309 747 3321 781
rect 3129 741 3321 747
rect -3377 697 -3331 709
rect -3377 121 -3371 697
rect -3337 121 -3331 697
rect -3377 109 -3331 121
rect -3119 697 -3073 709
rect -3119 121 -3113 697
rect -3079 121 -3073 697
rect -3119 109 -3073 121
rect -2861 697 -2815 709
rect -2861 121 -2855 697
rect -2821 121 -2815 697
rect -2861 109 -2815 121
rect -2603 697 -2557 709
rect -2603 121 -2597 697
rect -2563 121 -2557 697
rect -2603 109 -2557 121
rect -2345 697 -2299 709
rect -2345 121 -2339 697
rect -2305 121 -2299 697
rect -2345 109 -2299 121
rect -2087 697 -2041 709
rect -2087 121 -2081 697
rect -2047 121 -2041 697
rect -2087 109 -2041 121
rect -1829 697 -1783 709
rect -1829 121 -1823 697
rect -1789 121 -1783 697
rect -1829 109 -1783 121
rect -1571 697 -1525 709
rect -1571 121 -1565 697
rect -1531 121 -1525 697
rect -1571 109 -1525 121
rect -1313 697 -1267 709
rect -1313 121 -1307 697
rect -1273 121 -1267 697
rect -1313 109 -1267 121
rect -1055 697 -1009 709
rect -1055 121 -1049 697
rect -1015 121 -1009 697
rect -1055 109 -1009 121
rect -797 697 -751 709
rect -797 121 -791 697
rect -757 121 -751 697
rect -797 109 -751 121
rect -539 697 -493 709
rect -539 121 -533 697
rect -499 121 -493 697
rect -539 109 -493 121
rect -281 697 -235 709
rect -281 121 -275 697
rect -241 121 -235 697
rect -281 109 -235 121
rect -23 697 23 709
rect -23 121 -17 697
rect 17 121 23 697
rect -23 109 23 121
rect 235 697 281 709
rect 235 121 241 697
rect 275 121 281 697
rect 235 109 281 121
rect 493 697 539 709
rect 493 121 499 697
rect 533 121 539 697
rect 493 109 539 121
rect 751 697 797 709
rect 751 121 757 697
rect 791 121 797 697
rect 751 109 797 121
rect 1009 697 1055 709
rect 1009 121 1015 697
rect 1049 121 1055 697
rect 1009 109 1055 121
rect 1267 697 1313 709
rect 1267 121 1273 697
rect 1307 121 1313 697
rect 1267 109 1313 121
rect 1525 697 1571 709
rect 1525 121 1531 697
rect 1565 121 1571 697
rect 1525 109 1571 121
rect 1783 697 1829 709
rect 1783 121 1789 697
rect 1823 121 1829 697
rect 1783 109 1829 121
rect 2041 697 2087 709
rect 2041 121 2047 697
rect 2081 121 2087 697
rect 2041 109 2087 121
rect 2299 697 2345 709
rect 2299 121 2305 697
rect 2339 121 2345 697
rect 2299 109 2345 121
rect 2557 697 2603 709
rect 2557 121 2563 697
rect 2597 121 2603 697
rect 2557 109 2603 121
rect 2815 697 2861 709
rect 2815 121 2821 697
rect 2855 121 2861 697
rect 2815 109 2861 121
rect 3073 697 3119 709
rect 3073 121 3079 697
rect 3113 121 3119 697
rect 3073 109 3119 121
rect 3331 697 3377 709
rect 3331 121 3337 697
rect 3371 121 3377 697
rect 3331 109 3377 121
rect -3321 71 -3129 77
rect -3321 37 -3309 71
rect -3141 37 -3129 71
rect -3321 31 -3129 37
rect -3063 71 -2871 77
rect -3063 37 -3051 71
rect -2883 37 -2871 71
rect -3063 31 -2871 37
rect -2805 71 -2613 77
rect -2805 37 -2793 71
rect -2625 37 -2613 71
rect -2805 31 -2613 37
rect -2547 71 -2355 77
rect -2547 37 -2535 71
rect -2367 37 -2355 71
rect -2547 31 -2355 37
rect -2289 71 -2097 77
rect -2289 37 -2277 71
rect -2109 37 -2097 71
rect -2289 31 -2097 37
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect 2097 71 2289 77
rect 2097 37 2109 71
rect 2277 37 2289 71
rect 2097 31 2289 37
rect 2355 71 2547 77
rect 2355 37 2367 71
rect 2535 37 2547 71
rect 2355 31 2547 37
rect 2613 71 2805 77
rect 2613 37 2625 71
rect 2793 37 2805 71
rect 2613 31 2805 37
rect 2871 71 3063 77
rect 2871 37 2883 71
rect 3051 37 3063 71
rect 2871 31 3063 37
rect 3129 71 3321 77
rect 3129 37 3141 71
rect 3309 37 3321 71
rect 3129 31 3321 37
rect -3321 -37 -3129 -31
rect -3321 -71 -3309 -37
rect -3141 -71 -3129 -37
rect -3321 -77 -3129 -71
rect -3063 -37 -2871 -31
rect -3063 -71 -3051 -37
rect -2883 -71 -2871 -37
rect -3063 -77 -2871 -71
rect -2805 -37 -2613 -31
rect -2805 -71 -2793 -37
rect -2625 -71 -2613 -37
rect -2805 -77 -2613 -71
rect -2547 -37 -2355 -31
rect -2547 -71 -2535 -37
rect -2367 -71 -2355 -37
rect -2547 -77 -2355 -71
rect -2289 -37 -2097 -31
rect -2289 -71 -2277 -37
rect -2109 -71 -2097 -37
rect -2289 -77 -2097 -71
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect 2097 -37 2289 -31
rect 2097 -71 2109 -37
rect 2277 -71 2289 -37
rect 2097 -77 2289 -71
rect 2355 -37 2547 -31
rect 2355 -71 2367 -37
rect 2535 -71 2547 -37
rect 2355 -77 2547 -71
rect 2613 -37 2805 -31
rect 2613 -71 2625 -37
rect 2793 -71 2805 -37
rect 2613 -77 2805 -71
rect 2871 -37 3063 -31
rect 2871 -71 2883 -37
rect 3051 -71 3063 -37
rect 2871 -77 3063 -71
rect 3129 -37 3321 -31
rect 3129 -71 3141 -37
rect 3309 -71 3321 -37
rect 3129 -77 3321 -71
rect -3377 -121 -3331 -109
rect -3377 -697 -3371 -121
rect -3337 -697 -3331 -121
rect -3377 -709 -3331 -697
rect -3119 -121 -3073 -109
rect -3119 -697 -3113 -121
rect -3079 -697 -3073 -121
rect -3119 -709 -3073 -697
rect -2861 -121 -2815 -109
rect -2861 -697 -2855 -121
rect -2821 -697 -2815 -121
rect -2861 -709 -2815 -697
rect -2603 -121 -2557 -109
rect -2603 -697 -2597 -121
rect -2563 -697 -2557 -121
rect -2603 -709 -2557 -697
rect -2345 -121 -2299 -109
rect -2345 -697 -2339 -121
rect -2305 -697 -2299 -121
rect -2345 -709 -2299 -697
rect -2087 -121 -2041 -109
rect -2087 -697 -2081 -121
rect -2047 -697 -2041 -121
rect -2087 -709 -2041 -697
rect -1829 -121 -1783 -109
rect -1829 -697 -1823 -121
rect -1789 -697 -1783 -121
rect -1829 -709 -1783 -697
rect -1571 -121 -1525 -109
rect -1571 -697 -1565 -121
rect -1531 -697 -1525 -121
rect -1571 -709 -1525 -697
rect -1313 -121 -1267 -109
rect -1313 -697 -1307 -121
rect -1273 -697 -1267 -121
rect -1313 -709 -1267 -697
rect -1055 -121 -1009 -109
rect -1055 -697 -1049 -121
rect -1015 -697 -1009 -121
rect -1055 -709 -1009 -697
rect -797 -121 -751 -109
rect -797 -697 -791 -121
rect -757 -697 -751 -121
rect -797 -709 -751 -697
rect -539 -121 -493 -109
rect -539 -697 -533 -121
rect -499 -697 -493 -121
rect -539 -709 -493 -697
rect -281 -121 -235 -109
rect -281 -697 -275 -121
rect -241 -697 -235 -121
rect -281 -709 -235 -697
rect -23 -121 23 -109
rect -23 -697 -17 -121
rect 17 -697 23 -121
rect -23 -709 23 -697
rect 235 -121 281 -109
rect 235 -697 241 -121
rect 275 -697 281 -121
rect 235 -709 281 -697
rect 493 -121 539 -109
rect 493 -697 499 -121
rect 533 -697 539 -121
rect 493 -709 539 -697
rect 751 -121 797 -109
rect 751 -697 757 -121
rect 791 -697 797 -121
rect 751 -709 797 -697
rect 1009 -121 1055 -109
rect 1009 -697 1015 -121
rect 1049 -697 1055 -121
rect 1009 -709 1055 -697
rect 1267 -121 1313 -109
rect 1267 -697 1273 -121
rect 1307 -697 1313 -121
rect 1267 -709 1313 -697
rect 1525 -121 1571 -109
rect 1525 -697 1531 -121
rect 1565 -697 1571 -121
rect 1525 -709 1571 -697
rect 1783 -121 1829 -109
rect 1783 -697 1789 -121
rect 1823 -697 1829 -121
rect 1783 -709 1829 -697
rect 2041 -121 2087 -109
rect 2041 -697 2047 -121
rect 2081 -697 2087 -121
rect 2041 -709 2087 -697
rect 2299 -121 2345 -109
rect 2299 -697 2305 -121
rect 2339 -697 2345 -121
rect 2299 -709 2345 -697
rect 2557 -121 2603 -109
rect 2557 -697 2563 -121
rect 2597 -697 2603 -121
rect 2557 -709 2603 -697
rect 2815 -121 2861 -109
rect 2815 -697 2821 -121
rect 2855 -697 2861 -121
rect 2815 -709 2861 -697
rect 3073 -121 3119 -109
rect 3073 -697 3079 -121
rect 3113 -697 3119 -121
rect 3073 -709 3119 -697
rect 3331 -121 3377 -109
rect 3331 -697 3337 -121
rect 3371 -697 3377 -121
rect 3331 -709 3377 -697
rect -3321 -747 -3129 -741
rect -3321 -781 -3309 -747
rect -3141 -781 -3129 -747
rect -3321 -787 -3129 -781
rect -3063 -747 -2871 -741
rect -3063 -781 -3051 -747
rect -2883 -781 -2871 -747
rect -3063 -787 -2871 -781
rect -2805 -747 -2613 -741
rect -2805 -781 -2793 -747
rect -2625 -781 -2613 -747
rect -2805 -787 -2613 -781
rect -2547 -747 -2355 -741
rect -2547 -781 -2535 -747
rect -2367 -781 -2355 -747
rect -2547 -787 -2355 -781
rect -2289 -747 -2097 -741
rect -2289 -781 -2277 -747
rect -2109 -781 -2097 -747
rect -2289 -787 -2097 -781
rect -2031 -747 -1839 -741
rect -2031 -781 -2019 -747
rect -1851 -781 -1839 -747
rect -2031 -787 -1839 -781
rect -1773 -747 -1581 -741
rect -1773 -781 -1761 -747
rect -1593 -781 -1581 -747
rect -1773 -787 -1581 -781
rect -1515 -747 -1323 -741
rect -1515 -781 -1503 -747
rect -1335 -781 -1323 -747
rect -1515 -787 -1323 -781
rect -1257 -747 -1065 -741
rect -1257 -781 -1245 -747
rect -1077 -781 -1065 -747
rect -1257 -787 -1065 -781
rect -999 -747 -807 -741
rect -999 -781 -987 -747
rect -819 -781 -807 -747
rect -999 -787 -807 -781
rect -741 -747 -549 -741
rect -741 -781 -729 -747
rect -561 -781 -549 -747
rect -741 -787 -549 -781
rect -483 -747 -291 -741
rect -483 -781 -471 -747
rect -303 -781 -291 -747
rect -483 -787 -291 -781
rect -225 -747 -33 -741
rect -225 -781 -213 -747
rect -45 -781 -33 -747
rect -225 -787 -33 -781
rect 33 -747 225 -741
rect 33 -781 45 -747
rect 213 -781 225 -747
rect 33 -787 225 -781
rect 291 -747 483 -741
rect 291 -781 303 -747
rect 471 -781 483 -747
rect 291 -787 483 -781
rect 549 -747 741 -741
rect 549 -781 561 -747
rect 729 -781 741 -747
rect 549 -787 741 -781
rect 807 -747 999 -741
rect 807 -781 819 -747
rect 987 -781 999 -747
rect 807 -787 999 -781
rect 1065 -747 1257 -741
rect 1065 -781 1077 -747
rect 1245 -781 1257 -747
rect 1065 -787 1257 -781
rect 1323 -747 1515 -741
rect 1323 -781 1335 -747
rect 1503 -781 1515 -747
rect 1323 -787 1515 -781
rect 1581 -747 1773 -741
rect 1581 -781 1593 -747
rect 1761 -781 1773 -747
rect 1581 -787 1773 -781
rect 1839 -747 2031 -741
rect 1839 -781 1851 -747
rect 2019 -781 2031 -747
rect 1839 -787 2031 -781
rect 2097 -747 2289 -741
rect 2097 -781 2109 -747
rect 2277 -781 2289 -747
rect 2097 -787 2289 -781
rect 2355 -747 2547 -741
rect 2355 -781 2367 -747
rect 2535 -781 2547 -747
rect 2355 -787 2547 -781
rect 2613 -747 2805 -741
rect 2613 -781 2625 -747
rect 2793 -781 2805 -747
rect 2613 -787 2805 -781
rect 2871 -747 3063 -741
rect 2871 -781 2883 -747
rect 3051 -781 3063 -747
rect 2871 -787 3063 -781
rect 3129 -747 3321 -741
rect 3129 -781 3141 -747
rect 3309 -781 3321 -747
rect 3129 -787 3321 -781
<< properties >>
string FIXED_BBOX -3488 -902 3488 902
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3 l 1 m 2 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713300479
<< pwell >>
rect -4585 -1258 4585 1258
<< mvnmos >>
rect -4357 -1000 -4157 1000
rect -4099 -1000 -3899 1000
rect -3841 -1000 -3641 1000
rect -3583 -1000 -3383 1000
rect -3325 -1000 -3125 1000
rect -3067 -1000 -2867 1000
rect -2809 -1000 -2609 1000
rect -2551 -1000 -2351 1000
rect -2293 -1000 -2093 1000
rect -2035 -1000 -1835 1000
rect -1777 -1000 -1577 1000
rect -1519 -1000 -1319 1000
rect -1261 -1000 -1061 1000
rect -1003 -1000 -803 1000
rect -745 -1000 -545 1000
rect -487 -1000 -287 1000
rect -229 -1000 -29 1000
rect 29 -1000 229 1000
rect 287 -1000 487 1000
rect 545 -1000 745 1000
rect 803 -1000 1003 1000
rect 1061 -1000 1261 1000
rect 1319 -1000 1519 1000
rect 1577 -1000 1777 1000
rect 1835 -1000 2035 1000
rect 2093 -1000 2293 1000
rect 2351 -1000 2551 1000
rect 2609 -1000 2809 1000
rect 2867 -1000 3067 1000
rect 3125 -1000 3325 1000
rect 3383 -1000 3583 1000
rect 3641 -1000 3841 1000
rect 3899 -1000 4099 1000
rect 4157 -1000 4357 1000
<< mvndiff >>
rect -4415 988 -4357 1000
rect -4415 -988 -4403 988
rect -4369 -988 -4357 988
rect -4415 -1000 -4357 -988
rect -4157 988 -4099 1000
rect -4157 -988 -4145 988
rect -4111 -988 -4099 988
rect -4157 -1000 -4099 -988
rect -3899 988 -3841 1000
rect -3899 -988 -3887 988
rect -3853 -988 -3841 988
rect -3899 -1000 -3841 -988
rect -3641 988 -3583 1000
rect -3641 -988 -3629 988
rect -3595 -988 -3583 988
rect -3641 -1000 -3583 -988
rect -3383 988 -3325 1000
rect -3383 -988 -3371 988
rect -3337 -988 -3325 988
rect -3383 -1000 -3325 -988
rect -3125 988 -3067 1000
rect -3125 -988 -3113 988
rect -3079 -988 -3067 988
rect -3125 -1000 -3067 -988
rect -2867 988 -2809 1000
rect -2867 -988 -2855 988
rect -2821 -988 -2809 988
rect -2867 -1000 -2809 -988
rect -2609 988 -2551 1000
rect -2609 -988 -2597 988
rect -2563 -988 -2551 988
rect -2609 -1000 -2551 -988
rect -2351 988 -2293 1000
rect -2351 -988 -2339 988
rect -2305 -988 -2293 988
rect -2351 -1000 -2293 -988
rect -2093 988 -2035 1000
rect -2093 -988 -2081 988
rect -2047 -988 -2035 988
rect -2093 -1000 -2035 -988
rect -1835 988 -1777 1000
rect -1835 -988 -1823 988
rect -1789 -988 -1777 988
rect -1835 -1000 -1777 -988
rect -1577 988 -1519 1000
rect -1577 -988 -1565 988
rect -1531 -988 -1519 988
rect -1577 -1000 -1519 -988
rect -1319 988 -1261 1000
rect -1319 -988 -1307 988
rect -1273 -988 -1261 988
rect -1319 -1000 -1261 -988
rect -1061 988 -1003 1000
rect -1061 -988 -1049 988
rect -1015 -988 -1003 988
rect -1061 -1000 -1003 -988
rect -803 988 -745 1000
rect -803 -988 -791 988
rect -757 -988 -745 988
rect -803 -1000 -745 -988
rect -545 988 -487 1000
rect -545 -988 -533 988
rect -499 -988 -487 988
rect -545 -1000 -487 -988
rect -287 988 -229 1000
rect -287 -988 -275 988
rect -241 -988 -229 988
rect -287 -1000 -229 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 229 988 287 1000
rect 229 -988 241 988
rect 275 -988 287 988
rect 229 -1000 287 -988
rect 487 988 545 1000
rect 487 -988 499 988
rect 533 -988 545 988
rect 487 -1000 545 -988
rect 745 988 803 1000
rect 745 -988 757 988
rect 791 -988 803 988
rect 745 -1000 803 -988
rect 1003 988 1061 1000
rect 1003 -988 1015 988
rect 1049 -988 1061 988
rect 1003 -1000 1061 -988
rect 1261 988 1319 1000
rect 1261 -988 1273 988
rect 1307 -988 1319 988
rect 1261 -1000 1319 -988
rect 1519 988 1577 1000
rect 1519 -988 1531 988
rect 1565 -988 1577 988
rect 1519 -1000 1577 -988
rect 1777 988 1835 1000
rect 1777 -988 1789 988
rect 1823 -988 1835 988
rect 1777 -1000 1835 -988
rect 2035 988 2093 1000
rect 2035 -988 2047 988
rect 2081 -988 2093 988
rect 2035 -1000 2093 -988
rect 2293 988 2351 1000
rect 2293 -988 2305 988
rect 2339 -988 2351 988
rect 2293 -1000 2351 -988
rect 2551 988 2609 1000
rect 2551 -988 2563 988
rect 2597 -988 2609 988
rect 2551 -1000 2609 -988
rect 2809 988 2867 1000
rect 2809 -988 2821 988
rect 2855 -988 2867 988
rect 2809 -1000 2867 -988
rect 3067 988 3125 1000
rect 3067 -988 3079 988
rect 3113 -988 3125 988
rect 3067 -1000 3125 -988
rect 3325 988 3383 1000
rect 3325 -988 3337 988
rect 3371 -988 3383 988
rect 3325 -1000 3383 -988
rect 3583 988 3641 1000
rect 3583 -988 3595 988
rect 3629 -988 3641 988
rect 3583 -1000 3641 -988
rect 3841 988 3899 1000
rect 3841 -988 3853 988
rect 3887 -988 3899 988
rect 3841 -1000 3899 -988
rect 4099 988 4157 1000
rect 4099 -988 4111 988
rect 4145 -988 4157 988
rect 4099 -1000 4157 -988
rect 4357 988 4415 1000
rect 4357 -988 4369 988
rect 4403 -988 4415 988
rect 4357 -1000 4415 -988
<< mvndiffc >>
rect -4403 -988 -4369 988
rect -4145 -988 -4111 988
rect -3887 -988 -3853 988
rect -3629 -988 -3595 988
rect -3371 -988 -3337 988
rect -3113 -988 -3079 988
rect -2855 -988 -2821 988
rect -2597 -988 -2563 988
rect -2339 -988 -2305 988
rect -2081 -988 -2047 988
rect -1823 -988 -1789 988
rect -1565 -988 -1531 988
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect 1531 -988 1565 988
rect 1789 -988 1823 988
rect 2047 -988 2081 988
rect 2305 -988 2339 988
rect 2563 -988 2597 988
rect 2821 -988 2855 988
rect 3079 -988 3113 988
rect 3337 -988 3371 988
rect 3595 -988 3629 988
rect 3853 -988 3887 988
rect 4111 -988 4145 988
rect 4369 -988 4403 988
<< mvpsubdiff >>
rect -4549 1210 4549 1222
rect -4549 1176 -4441 1210
rect 4441 1176 4549 1210
rect -4549 1164 4549 1176
rect -4549 1114 -4491 1164
rect -4549 -1114 -4537 1114
rect -4503 -1114 -4491 1114
rect 4491 1114 4549 1164
rect -4549 -1164 -4491 -1114
rect 4491 -1114 4503 1114
rect 4537 -1114 4549 1114
rect 4491 -1164 4549 -1114
rect -4549 -1176 4549 -1164
rect -4549 -1210 -4441 -1176
rect 4441 -1210 4549 -1176
rect -4549 -1222 4549 -1210
<< mvpsubdiffcont >>
rect -4441 1176 4441 1210
rect -4537 -1114 -4503 1114
rect 4503 -1114 4537 1114
rect -4441 -1210 4441 -1176
<< poly >>
rect -4323 1072 -4191 1088
rect -4323 1055 -4307 1072
rect -4357 1038 -4307 1055
rect -4207 1055 -4191 1072
rect -4065 1072 -3933 1088
rect -4065 1055 -4049 1072
rect -4207 1038 -4157 1055
rect -4357 1000 -4157 1038
rect -4099 1038 -4049 1055
rect -3949 1055 -3933 1072
rect -3807 1072 -3675 1088
rect -3807 1055 -3791 1072
rect -3949 1038 -3899 1055
rect -4099 1000 -3899 1038
rect -3841 1038 -3791 1055
rect -3691 1055 -3675 1072
rect -3549 1072 -3417 1088
rect -3549 1055 -3533 1072
rect -3691 1038 -3641 1055
rect -3841 1000 -3641 1038
rect -3583 1038 -3533 1055
rect -3433 1055 -3417 1072
rect -3291 1072 -3159 1088
rect -3291 1055 -3275 1072
rect -3433 1038 -3383 1055
rect -3583 1000 -3383 1038
rect -3325 1038 -3275 1055
rect -3175 1055 -3159 1072
rect -3033 1072 -2901 1088
rect -3033 1055 -3017 1072
rect -3175 1038 -3125 1055
rect -3325 1000 -3125 1038
rect -3067 1038 -3017 1055
rect -2917 1055 -2901 1072
rect -2775 1072 -2643 1088
rect -2775 1055 -2759 1072
rect -2917 1038 -2867 1055
rect -3067 1000 -2867 1038
rect -2809 1038 -2759 1055
rect -2659 1055 -2643 1072
rect -2517 1072 -2385 1088
rect -2517 1055 -2501 1072
rect -2659 1038 -2609 1055
rect -2809 1000 -2609 1038
rect -2551 1038 -2501 1055
rect -2401 1055 -2385 1072
rect -2259 1072 -2127 1088
rect -2259 1055 -2243 1072
rect -2401 1038 -2351 1055
rect -2551 1000 -2351 1038
rect -2293 1038 -2243 1055
rect -2143 1055 -2127 1072
rect -2001 1072 -1869 1088
rect -2001 1055 -1985 1072
rect -2143 1038 -2093 1055
rect -2293 1000 -2093 1038
rect -2035 1038 -1985 1055
rect -1885 1055 -1869 1072
rect -1743 1072 -1611 1088
rect -1743 1055 -1727 1072
rect -1885 1038 -1835 1055
rect -2035 1000 -1835 1038
rect -1777 1038 -1727 1055
rect -1627 1055 -1611 1072
rect -1485 1072 -1353 1088
rect -1485 1055 -1469 1072
rect -1627 1038 -1577 1055
rect -1777 1000 -1577 1038
rect -1519 1038 -1469 1055
rect -1369 1055 -1353 1072
rect -1227 1072 -1095 1088
rect -1227 1055 -1211 1072
rect -1369 1038 -1319 1055
rect -1519 1000 -1319 1038
rect -1261 1038 -1211 1055
rect -1111 1055 -1095 1072
rect -969 1072 -837 1088
rect -969 1055 -953 1072
rect -1111 1038 -1061 1055
rect -1261 1000 -1061 1038
rect -1003 1038 -953 1055
rect -853 1055 -837 1072
rect -711 1072 -579 1088
rect -711 1055 -695 1072
rect -853 1038 -803 1055
rect -1003 1000 -803 1038
rect -745 1038 -695 1055
rect -595 1055 -579 1072
rect -453 1072 -321 1088
rect -453 1055 -437 1072
rect -595 1038 -545 1055
rect -745 1000 -545 1038
rect -487 1038 -437 1055
rect -337 1055 -321 1072
rect -195 1072 -63 1088
rect -195 1055 -179 1072
rect -337 1038 -287 1055
rect -487 1000 -287 1038
rect -229 1038 -179 1055
rect -79 1055 -63 1072
rect 63 1072 195 1088
rect 63 1055 79 1072
rect -79 1038 -29 1055
rect -229 1000 -29 1038
rect 29 1038 79 1055
rect 179 1055 195 1072
rect 321 1072 453 1088
rect 321 1055 337 1072
rect 179 1038 229 1055
rect 29 1000 229 1038
rect 287 1038 337 1055
rect 437 1055 453 1072
rect 579 1072 711 1088
rect 579 1055 595 1072
rect 437 1038 487 1055
rect 287 1000 487 1038
rect 545 1038 595 1055
rect 695 1055 711 1072
rect 837 1072 969 1088
rect 837 1055 853 1072
rect 695 1038 745 1055
rect 545 1000 745 1038
rect 803 1038 853 1055
rect 953 1055 969 1072
rect 1095 1072 1227 1088
rect 1095 1055 1111 1072
rect 953 1038 1003 1055
rect 803 1000 1003 1038
rect 1061 1038 1111 1055
rect 1211 1055 1227 1072
rect 1353 1072 1485 1088
rect 1353 1055 1369 1072
rect 1211 1038 1261 1055
rect 1061 1000 1261 1038
rect 1319 1038 1369 1055
rect 1469 1055 1485 1072
rect 1611 1072 1743 1088
rect 1611 1055 1627 1072
rect 1469 1038 1519 1055
rect 1319 1000 1519 1038
rect 1577 1038 1627 1055
rect 1727 1055 1743 1072
rect 1869 1072 2001 1088
rect 1869 1055 1885 1072
rect 1727 1038 1777 1055
rect 1577 1000 1777 1038
rect 1835 1038 1885 1055
rect 1985 1055 2001 1072
rect 2127 1072 2259 1088
rect 2127 1055 2143 1072
rect 1985 1038 2035 1055
rect 1835 1000 2035 1038
rect 2093 1038 2143 1055
rect 2243 1055 2259 1072
rect 2385 1072 2517 1088
rect 2385 1055 2401 1072
rect 2243 1038 2293 1055
rect 2093 1000 2293 1038
rect 2351 1038 2401 1055
rect 2501 1055 2517 1072
rect 2643 1072 2775 1088
rect 2643 1055 2659 1072
rect 2501 1038 2551 1055
rect 2351 1000 2551 1038
rect 2609 1038 2659 1055
rect 2759 1055 2775 1072
rect 2901 1072 3033 1088
rect 2901 1055 2917 1072
rect 2759 1038 2809 1055
rect 2609 1000 2809 1038
rect 2867 1038 2917 1055
rect 3017 1055 3033 1072
rect 3159 1072 3291 1088
rect 3159 1055 3175 1072
rect 3017 1038 3067 1055
rect 2867 1000 3067 1038
rect 3125 1038 3175 1055
rect 3275 1055 3291 1072
rect 3417 1072 3549 1088
rect 3417 1055 3433 1072
rect 3275 1038 3325 1055
rect 3125 1000 3325 1038
rect 3383 1038 3433 1055
rect 3533 1055 3549 1072
rect 3675 1072 3807 1088
rect 3675 1055 3691 1072
rect 3533 1038 3583 1055
rect 3383 1000 3583 1038
rect 3641 1038 3691 1055
rect 3791 1055 3807 1072
rect 3933 1072 4065 1088
rect 3933 1055 3949 1072
rect 3791 1038 3841 1055
rect 3641 1000 3841 1038
rect 3899 1038 3949 1055
rect 4049 1055 4065 1072
rect 4191 1072 4323 1088
rect 4191 1055 4207 1072
rect 4049 1038 4099 1055
rect 3899 1000 4099 1038
rect 4157 1038 4207 1055
rect 4307 1055 4323 1072
rect 4307 1038 4357 1055
rect 4157 1000 4357 1038
rect -4357 -1038 -4157 -1000
rect -4357 -1055 -4307 -1038
rect -4323 -1072 -4307 -1055
rect -4207 -1055 -4157 -1038
rect -4099 -1038 -3899 -1000
rect -4099 -1055 -4049 -1038
rect -4207 -1072 -4191 -1055
rect -4323 -1088 -4191 -1072
rect -4065 -1072 -4049 -1055
rect -3949 -1055 -3899 -1038
rect -3841 -1038 -3641 -1000
rect -3841 -1055 -3791 -1038
rect -3949 -1072 -3933 -1055
rect -4065 -1088 -3933 -1072
rect -3807 -1072 -3791 -1055
rect -3691 -1055 -3641 -1038
rect -3583 -1038 -3383 -1000
rect -3583 -1055 -3533 -1038
rect -3691 -1072 -3675 -1055
rect -3807 -1088 -3675 -1072
rect -3549 -1072 -3533 -1055
rect -3433 -1055 -3383 -1038
rect -3325 -1038 -3125 -1000
rect -3325 -1055 -3275 -1038
rect -3433 -1072 -3417 -1055
rect -3549 -1088 -3417 -1072
rect -3291 -1072 -3275 -1055
rect -3175 -1055 -3125 -1038
rect -3067 -1038 -2867 -1000
rect -3067 -1055 -3017 -1038
rect -3175 -1072 -3159 -1055
rect -3291 -1088 -3159 -1072
rect -3033 -1072 -3017 -1055
rect -2917 -1055 -2867 -1038
rect -2809 -1038 -2609 -1000
rect -2809 -1055 -2759 -1038
rect -2917 -1072 -2901 -1055
rect -3033 -1088 -2901 -1072
rect -2775 -1072 -2759 -1055
rect -2659 -1055 -2609 -1038
rect -2551 -1038 -2351 -1000
rect -2551 -1055 -2501 -1038
rect -2659 -1072 -2643 -1055
rect -2775 -1088 -2643 -1072
rect -2517 -1072 -2501 -1055
rect -2401 -1055 -2351 -1038
rect -2293 -1038 -2093 -1000
rect -2293 -1055 -2243 -1038
rect -2401 -1072 -2385 -1055
rect -2517 -1088 -2385 -1072
rect -2259 -1072 -2243 -1055
rect -2143 -1055 -2093 -1038
rect -2035 -1038 -1835 -1000
rect -2035 -1055 -1985 -1038
rect -2143 -1072 -2127 -1055
rect -2259 -1088 -2127 -1072
rect -2001 -1072 -1985 -1055
rect -1885 -1055 -1835 -1038
rect -1777 -1038 -1577 -1000
rect -1777 -1055 -1727 -1038
rect -1885 -1072 -1869 -1055
rect -2001 -1088 -1869 -1072
rect -1743 -1072 -1727 -1055
rect -1627 -1055 -1577 -1038
rect -1519 -1038 -1319 -1000
rect -1519 -1055 -1469 -1038
rect -1627 -1072 -1611 -1055
rect -1743 -1088 -1611 -1072
rect -1485 -1072 -1469 -1055
rect -1369 -1055 -1319 -1038
rect -1261 -1038 -1061 -1000
rect -1261 -1055 -1211 -1038
rect -1369 -1072 -1353 -1055
rect -1485 -1088 -1353 -1072
rect -1227 -1072 -1211 -1055
rect -1111 -1055 -1061 -1038
rect -1003 -1038 -803 -1000
rect -1003 -1055 -953 -1038
rect -1111 -1072 -1095 -1055
rect -1227 -1088 -1095 -1072
rect -969 -1072 -953 -1055
rect -853 -1055 -803 -1038
rect -745 -1038 -545 -1000
rect -745 -1055 -695 -1038
rect -853 -1072 -837 -1055
rect -969 -1088 -837 -1072
rect -711 -1072 -695 -1055
rect -595 -1055 -545 -1038
rect -487 -1038 -287 -1000
rect -487 -1055 -437 -1038
rect -595 -1072 -579 -1055
rect -711 -1088 -579 -1072
rect -453 -1072 -437 -1055
rect -337 -1055 -287 -1038
rect -229 -1038 -29 -1000
rect -229 -1055 -179 -1038
rect -337 -1072 -321 -1055
rect -453 -1088 -321 -1072
rect -195 -1072 -179 -1055
rect -79 -1055 -29 -1038
rect 29 -1038 229 -1000
rect 29 -1055 79 -1038
rect -79 -1072 -63 -1055
rect -195 -1088 -63 -1072
rect 63 -1072 79 -1055
rect 179 -1055 229 -1038
rect 287 -1038 487 -1000
rect 287 -1055 337 -1038
rect 179 -1072 195 -1055
rect 63 -1088 195 -1072
rect 321 -1072 337 -1055
rect 437 -1055 487 -1038
rect 545 -1038 745 -1000
rect 545 -1055 595 -1038
rect 437 -1072 453 -1055
rect 321 -1088 453 -1072
rect 579 -1072 595 -1055
rect 695 -1055 745 -1038
rect 803 -1038 1003 -1000
rect 803 -1055 853 -1038
rect 695 -1072 711 -1055
rect 579 -1088 711 -1072
rect 837 -1072 853 -1055
rect 953 -1055 1003 -1038
rect 1061 -1038 1261 -1000
rect 1061 -1055 1111 -1038
rect 953 -1072 969 -1055
rect 837 -1088 969 -1072
rect 1095 -1072 1111 -1055
rect 1211 -1055 1261 -1038
rect 1319 -1038 1519 -1000
rect 1319 -1055 1369 -1038
rect 1211 -1072 1227 -1055
rect 1095 -1088 1227 -1072
rect 1353 -1072 1369 -1055
rect 1469 -1055 1519 -1038
rect 1577 -1038 1777 -1000
rect 1577 -1055 1627 -1038
rect 1469 -1072 1485 -1055
rect 1353 -1088 1485 -1072
rect 1611 -1072 1627 -1055
rect 1727 -1055 1777 -1038
rect 1835 -1038 2035 -1000
rect 1835 -1055 1885 -1038
rect 1727 -1072 1743 -1055
rect 1611 -1088 1743 -1072
rect 1869 -1072 1885 -1055
rect 1985 -1055 2035 -1038
rect 2093 -1038 2293 -1000
rect 2093 -1055 2143 -1038
rect 1985 -1072 2001 -1055
rect 1869 -1088 2001 -1072
rect 2127 -1072 2143 -1055
rect 2243 -1055 2293 -1038
rect 2351 -1038 2551 -1000
rect 2351 -1055 2401 -1038
rect 2243 -1072 2259 -1055
rect 2127 -1088 2259 -1072
rect 2385 -1072 2401 -1055
rect 2501 -1055 2551 -1038
rect 2609 -1038 2809 -1000
rect 2609 -1055 2659 -1038
rect 2501 -1072 2517 -1055
rect 2385 -1088 2517 -1072
rect 2643 -1072 2659 -1055
rect 2759 -1055 2809 -1038
rect 2867 -1038 3067 -1000
rect 2867 -1055 2917 -1038
rect 2759 -1072 2775 -1055
rect 2643 -1088 2775 -1072
rect 2901 -1072 2917 -1055
rect 3017 -1055 3067 -1038
rect 3125 -1038 3325 -1000
rect 3125 -1055 3175 -1038
rect 3017 -1072 3033 -1055
rect 2901 -1088 3033 -1072
rect 3159 -1072 3175 -1055
rect 3275 -1055 3325 -1038
rect 3383 -1038 3583 -1000
rect 3383 -1055 3433 -1038
rect 3275 -1072 3291 -1055
rect 3159 -1088 3291 -1072
rect 3417 -1072 3433 -1055
rect 3533 -1055 3583 -1038
rect 3641 -1038 3841 -1000
rect 3641 -1055 3691 -1038
rect 3533 -1072 3549 -1055
rect 3417 -1088 3549 -1072
rect 3675 -1072 3691 -1055
rect 3791 -1055 3841 -1038
rect 3899 -1038 4099 -1000
rect 3899 -1055 3949 -1038
rect 3791 -1072 3807 -1055
rect 3675 -1088 3807 -1072
rect 3933 -1072 3949 -1055
rect 4049 -1055 4099 -1038
rect 4157 -1038 4357 -1000
rect 4157 -1055 4207 -1038
rect 4049 -1072 4065 -1055
rect 3933 -1088 4065 -1072
rect 4191 -1072 4207 -1055
rect 4307 -1055 4357 -1038
rect 4307 -1072 4323 -1055
rect 4191 -1088 4323 -1072
<< polycont >>
rect -4307 1038 -4207 1072
rect -4049 1038 -3949 1072
rect -3791 1038 -3691 1072
rect -3533 1038 -3433 1072
rect -3275 1038 -3175 1072
rect -3017 1038 -2917 1072
rect -2759 1038 -2659 1072
rect -2501 1038 -2401 1072
rect -2243 1038 -2143 1072
rect -1985 1038 -1885 1072
rect -1727 1038 -1627 1072
rect -1469 1038 -1369 1072
rect -1211 1038 -1111 1072
rect -953 1038 -853 1072
rect -695 1038 -595 1072
rect -437 1038 -337 1072
rect -179 1038 -79 1072
rect 79 1038 179 1072
rect 337 1038 437 1072
rect 595 1038 695 1072
rect 853 1038 953 1072
rect 1111 1038 1211 1072
rect 1369 1038 1469 1072
rect 1627 1038 1727 1072
rect 1885 1038 1985 1072
rect 2143 1038 2243 1072
rect 2401 1038 2501 1072
rect 2659 1038 2759 1072
rect 2917 1038 3017 1072
rect 3175 1038 3275 1072
rect 3433 1038 3533 1072
rect 3691 1038 3791 1072
rect 3949 1038 4049 1072
rect 4207 1038 4307 1072
rect -4307 -1072 -4207 -1038
rect -4049 -1072 -3949 -1038
rect -3791 -1072 -3691 -1038
rect -3533 -1072 -3433 -1038
rect -3275 -1072 -3175 -1038
rect -3017 -1072 -2917 -1038
rect -2759 -1072 -2659 -1038
rect -2501 -1072 -2401 -1038
rect -2243 -1072 -2143 -1038
rect -1985 -1072 -1885 -1038
rect -1727 -1072 -1627 -1038
rect -1469 -1072 -1369 -1038
rect -1211 -1072 -1111 -1038
rect -953 -1072 -853 -1038
rect -695 -1072 -595 -1038
rect -437 -1072 -337 -1038
rect -179 -1072 -79 -1038
rect 79 -1072 179 -1038
rect 337 -1072 437 -1038
rect 595 -1072 695 -1038
rect 853 -1072 953 -1038
rect 1111 -1072 1211 -1038
rect 1369 -1072 1469 -1038
rect 1627 -1072 1727 -1038
rect 1885 -1072 1985 -1038
rect 2143 -1072 2243 -1038
rect 2401 -1072 2501 -1038
rect 2659 -1072 2759 -1038
rect 2917 -1072 3017 -1038
rect 3175 -1072 3275 -1038
rect 3433 -1072 3533 -1038
rect 3691 -1072 3791 -1038
rect 3949 -1072 4049 -1038
rect 4207 -1072 4307 -1038
<< locali >>
rect -4537 1176 -4441 1210
rect 4441 1176 4537 1210
rect -4537 1114 -4503 1176
rect 4503 1114 4537 1176
rect -4323 1038 -4307 1072
rect -4207 1038 -4191 1072
rect -4065 1038 -4049 1072
rect -3949 1038 -3933 1072
rect -3807 1038 -3791 1072
rect -3691 1038 -3675 1072
rect -3549 1038 -3533 1072
rect -3433 1038 -3417 1072
rect -3291 1038 -3275 1072
rect -3175 1038 -3159 1072
rect -3033 1038 -3017 1072
rect -2917 1038 -2901 1072
rect -2775 1038 -2759 1072
rect -2659 1038 -2643 1072
rect -2517 1038 -2501 1072
rect -2401 1038 -2385 1072
rect -2259 1038 -2243 1072
rect -2143 1038 -2127 1072
rect -2001 1038 -1985 1072
rect -1885 1038 -1869 1072
rect -1743 1038 -1727 1072
rect -1627 1038 -1611 1072
rect -1485 1038 -1469 1072
rect -1369 1038 -1353 1072
rect -1227 1038 -1211 1072
rect -1111 1038 -1095 1072
rect -969 1038 -953 1072
rect -853 1038 -837 1072
rect -711 1038 -695 1072
rect -595 1038 -579 1072
rect -453 1038 -437 1072
rect -337 1038 -321 1072
rect -195 1038 -179 1072
rect -79 1038 -63 1072
rect 63 1038 79 1072
rect 179 1038 195 1072
rect 321 1038 337 1072
rect 437 1038 453 1072
rect 579 1038 595 1072
rect 695 1038 711 1072
rect 837 1038 853 1072
rect 953 1038 969 1072
rect 1095 1038 1111 1072
rect 1211 1038 1227 1072
rect 1353 1038 1369 1072
rect 1469 1038 1485 1072
rect 1611 1038 1627 1072
rect 1727 1038 1743 1072
rect 1869 1038 1885 1072
rect 1985 1038 2001 1072
rect 2127 1038 2143 1072
rect 2243 1038 2259 1072
rect 2385 1038 2401 1072
rect 2501 1038 2517 1072
rect 2643 1038 2659 1072
rect 2759 1038 2775 1072
rect 2901 1038 2917 1072
rect 3017 1038 3033 1072
rect 3159 1038 3175 1072
rect 3275 1038 3291 1072
rect 3417 1038 3433 1072
rect 3533 1038 3549 1072
rect 3675 1038 3691 1072
rect 3791 1038 3807 1072
rect 3933 1038 3949 1072
rect 4049 1038 4065 1072
rect 4191 1038 4207 1072
rect 4307 1038 4323 1072
rect -4403 988 -4369 1004
rect -4403 -1004 -4369 -988
rect -4145 988 -4111 1004
rect -4145 -1004 -4111 -988
rect -3887 988 -3853 1004
rect -3887 -1004 -3853 -988
rect -3629 988 -3595 1004
rect -3629 -1004 -3595 -988
rect -3371 988 -3337 1004
rect -3371 -1004 -3337 -988
rect -3113 988 -3079 1004
rect -3113 -1004 -3079 -988
rect -2855 988 -2821 1004
rect -2855 -1004 -2821 -988
rect -2597 988 -2563 1004
rect -2597 -1004 -2563 -988
rect -2339 988 -2305 1004
rect -2339 -1004 -2305 -988
rect -2081 988 -2047 1004
rect -2081 -1004 -2047 -988
rect -1823 988 -1789 1004
rect -1823 -1004 -1789 -988
rect -1565 988 -1531 1004
rect -1565 -1004 -1531 -988
rect -1307 988 -1273 1004
rect -1307 -1004 -1273 -988
rect -1049 988 -1015 1004
rect -1049 -1004 -1015 -988
rect -791 988 -757 1004
rect -791 -1004 -757 -988
rect -533 988 -499 1004
rect -533 -1004 -499 -988
rect -275 988 -241 1004
rect -275 -1004 -241 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 241 988 275 1004
rect 241 -1004 275 -988
rect 499 988 533 1004
rect 499 -1004 533 -988
rect 757 988 791 1004
rect 757 -1004 791 -988
rect 1015 988 1049 1004
rect 1015 -1004 1049 -988
rect 1273 988 1307 1004
rect 1273 -1004 1307 -988
rect 1531 988 1565 1004
rect 1531 -1004 1565 -988
rect 1789 988 1823 1004
rect 1789 -1004 1823 -988
rect 2047 988 2081 1004
rect 2047 -1004 2081 -988
rect 2305 988 2339 1004
rect 2305 -1004 2339 -988
rect 2563 988 2597 1004
rect 2563 -1004 2597 -988
rect 2821 988 2855 1004
rect 2821 -1004 2855 -988
rect 3079 988 3113 1004
rect 3079 -1004 3113 -988
rect 3337 988 3371 1004
rect 3337 -1004 3371 -988
rect 3595 988 3629 1004
rect 3595 -1004 3629 -988
rect 3853 988 3887 1004
rect 3853 -1004 3887 -988
rect 4111 988 4145 1004
rect 4111 -1004 4145 -988
rect 4369 988 4403 1004
rect 4369 -1004 4403 -988
rect -4323 -1072 -4307 -1038
rect -4207 -1072 -4191 -1038
rect -4065 -1072 -4049 -1038
rect -3949 -1072 -3933 -1038
rect -3807 -1072 -3791 -1038
rect -3691 -1072 -3675 -1038
rect -3549 -1072 -3533 -1038
rect -3433 -1072 -3417 -1038
rect -3291 -1072 -3275 -1038
rect -3175 -1072 -3159 -1038
rect -3033 -1072 -3017 -1038
rect -2917 -1072 -2901 -1038
rect -2775 -1072 -2759 -1038
rect -2659 -1072 -2643 -1038
rect -2517 -1072 -2501 -1038
rect -2401 -1072 -2385 -1038
rect -2259 -1072 -2243 -1038
rect -2143 -1072 -2127 -1038
rect -2001 -1072 -1985 -1038
rect -1885 -1072 -1869 -1038
rect -1743 -1072 -1727 -1038
rect -1627 -1072 -1611 -1038
rect -1485 -1072 -1469 -1038
rect -1369 -1072 -1353 -1038
rect -1227 -1072 -1211 -1038
rect -1111 -1072 -1095 -1038
rect -969 -1072 -953 -1038
rect -853 -1072 -837 -1038
rect -711 -1072 -695 -1038
rect -595 -1072 -579 -1038
rect -453 -1072 -437 -1038
rect -337 -1072 -321 -1038
rect -195 -1072 -179 -1038
rect -79 -1072 -63 -1038
rect 63 -1072 79 -1038
rect 179 -1072 195 -1038
rect 321 -1072 337 -1038
rect 437 -1072 453 -1038
rect 579 -1072 595 -1038
rect 695 -1072 711 -1038
rect 837 -1072 853 -1038
rect 953 -1072 969 -1038
rect 1095 -1072 1111 -1038
rect 1211 -1072 1227 -1038
rect 1353 -1072 1369 -1038
rect 1469 -1072 1485 -1038
rect 1611 -1072 1627 -1038
rect 1727 -1072 1743 -1038
rect 1869 -1072 1885 -1038
rect 1985 -1072 2001 -1038
rect 2127 -1072 2143 -1038
rect 2243 -1072 2259 -1038
rect 2385 -1072 2401 -1038
rect 2501 -1072 2517 -1038
rect 2643 -1072 2659 -1038
rect 2759 -1072 2775 -1038
rect 2901 -1072 2917 -1038
rect 3017 -1072 3033 -1038
rect 3159 -1072 3175 -1038
rect 3275 -1072 3291 -1038
rect 3417 -1072 3433 -1038
rect 3533 -1072 3549 -1038
rect 3675 -1072 3691 -1038
rect 3791 -1072 3807 -1038
rect 3933 -1072 3949 -1038
rect 4049 -1072 4065 -1038
rect 4191 -1072 4207 -1038
rect 4307 -1072 4323 -1038
rect -4537 -1176 -4503 -1114
rect 4503 -1176 4537 -1114
rect -4537 -1210 -4441 -1176
rect 4441 -1210 4537 -1176
<< viali >>
rect -4307 1038 -4207 1072
rect -4049 1038 -3949 1072
rect -3791 1038 -3691 1072
rect -3533 1038 -3433 1072
rect -3275 1038 -3175 1072
rect -3017 1038 -2917 1072
rect -2759 1038 -2659 1072
rect -2501 1038 -2401 1072
rect -2243 1038 -2143 1072
rect -1985 1038 -1885 1072
rect -1727 1038 -1627 1072
rect -1469 1038 -1369 1072
rect -1211 1038 -1111 1072
rect -953 1038 -853 1072
rect -695 1038 -595 1072
rect -437 1038 -337 1072
rect -179 1038 -79 1072
rect 79 1038 179 1072
rect 337 1038 437 1072
rect 595 1038 695 1072
rect 853 1038 953 1072
rect 1111 1038 1211 1072
rect 1369 1038 1469 1072
rect 1627 1038 1727 1072
rect 1885 1038 1985 1072
rect 2143 1038 2243 1072
rect 2401 1038 2501 1072
rect 2659 1038 2759 1072
rect 2917 1038 3017 1072
rect 3175 1038 3275 1072
rect 3433 1038 3533 1072
rect 3691 1038 3791 1072
rect 3949 1038 4049 1072
rect 4207 1038 4307 1072
rect -4403 -988 -4369 988
rect -4145 -988 -4111 988
rect -3887 -988 -3853 988
rect -3629 -988 -3595 988
rect -3371 -988 -3337 988
rect -3113 -988 -3079 988
rect -2855 -988 -2821 988
rect -2597 -988 -2563 988
rect -2339 -988 -2305 988
rect -2081 -988 -2047 988
rect -1823 -988 -1789 988
rect -1565 -988 -1531 988
rect -1307 -988 -1273 988
rect -1049 -988 -1015 988
rect -791 -988 -757 988
rect -533 -988 -499 988
rect -275 -988 -241 988
rect -17 -988 17 988
rect 241 -988 275 988
rect 499 -988 533 988
rect 757 -988 791 988
rect 1015 -988 1049 988
rect 1273 -988 1307 988
rect 1531 -988 1565 988
rect 1789 -988 1823 988
rect 2047 -988 2081 988
rect 2305 -988 2339 988
rect 2563 -988 2597 988
rect 2821 -988 2855 988
rect 3079 -988 3113 988
rect 3337 -988 3371 988
rect 3595 -988 3629 988
rect 3853 -988 3887 988
rect 4111 -988 4145 988
rect 4369 -988 4403 988
rect -4307 -1072 -4207 -1038
rect -4049 -1072 -3949 -1038
rect -3791 -1072 -3691 -1038
rect -3533 -1072 -3433 -1038
rect -3275 -1072 -3175 -1038
rect -3017 -1072 -2917 -1038
rect -2759 -1072 -2659 -1038
rect -2501 -1072 -2401 -1038
rect -2243 -1072 -2143 -1038
rect -1985 -1072 -1885 -1038
rect -1727 -1072 -1627 -1038
rect -1469 -1072 -1369 -1038
rect -1211 -1072 -1111 -1038
rect -953 -1072 -853 -1038
rect -695 -1072 -595 -1038
rect -437 -1072 -337 -1038
rect -179 -1072 -79 -1038
rect 79 -1072 179 -1038
rect 337 -1072 437 -1038
rect 595 -1072 695 -1038
rect 853 -1072 953 -1038
rect 1111 -1072 1211 -1038
rect 1369 -1072 1469 -1038
rect 1627 -1072 1727 -1038
rect 1885 -1072 1985 -1038
rect 2143 -1072 2243 -1038
rect 2401 -1072 2501 -1038
rect 2659 -1072 2759 -1038
rect 2917 -1072 3017 -1038
rect 3175 -1072 3275 -1038
rect 3433 -1072 3533 -1038
rect 3691 -1072 3791 -1038
rect 3949 -1072 4049 -1038
rect 4207 -1072 4307 -1038
<< metal1 >>
rect -4319 1072 -4195 1078
rect -4319 1038 -4307 1072
rect -4207 1038 -4195 1072
rect -4319 1032 -4195 1038
rect -4061 1072 -3937 1078
rect -4061 1038 -4049 1072
rect -3949 1038 -3937 1072
rect -4061 1032 -3937 1038
rect -3803 1072 -3679 1078
rect -3803 1038 -3791 1072
rect -3691 1038 -3679 1072
rect -3803 1032 -3679 1038
rect -3545 1072 -3421 1078
rect -3545 1038 -3533 1072
rect -3433 1038 -3421 1072
rect -3545 1032 -3421 1038
rect -3287 1072 -3163 1078
rect -3287 1038 -3275 1072
rect -3175 1038 -3163 1072
rect -3287 1032 -3163 1038
rect -3029 1072 -2905 1078
rect -3029 1038 -3017 1072
rect -2917 1038 -2905 1072
rect -3029 1032 -2905 1038
rect -2771 1072 -2647 1078
rect -2771 1038 -2759 1072
rect -2659 1038 -2647 1072
rect -2771 1032 -2647 1038
rect -2513 1072 -2389 1078
rect -2513 1038 -2501 1072
rect -2401 1038 -2389 1072
rect -2513 1032 -2389 1038
rect -2255 1072 -2131 1078
rect -2255 1038 -2243 1072
rect -2143 1038 -2131 1072
rect -2255 1032 -2131 1038
rect -1997 1072 -1873 1078
rect -1997 1038 -1985 1072
rect -1885 1038 -1873 1072
rect -1997 1032 -1873 1038
rect -1739 1072 -1615 1078
rect -1739 1038 -1727 1072
rect -1627 1038 -1615 1072
rect -1739 1032 -1615 1038
rect -1481 1072 -1357 1078
rect -1481 1038 -1469 1072
rect -1369 1038 -1357 1072
rect -1481 1032 -1357 1038
rect -1223 1072 -1099 1078
rect -1223 1038 -1211 1072
rect -1111 1038 -1099 1072
rect -1223 1032 -1099 1038
rect -965 1072 -841 1078
rect -965 1038 -953 1072
rect -853 1038 -841 1072
rect -965 1032 -841 1038
rect -707 1072 -583 1078
rect -707 1038 -695 1072
rect -595 1038 -583 1072
rect -707 1032 -583 1038
rect -449 1072 -325 1078
rect -449 1038 -437 1072
rect -337 1038 -325 1072
rect -449 1032 -325 1038
rect -191 1072 -67 1078
rect -191 1038 -179 1072
rect -79 1038 -67 1072
rect -191 1032 -67 1038
rect 67 1072 191 1078
rect 67 1038 79 1072
rect 179 1038 191 1072
rect 67 1032 191 1038
rect 325 1072 449 1078
rect 325 1038 337 1072
rect 437 1038 449 1072
rect 325 1032 449 1038
rect 583 1072 707 1078
rect 583 1038 595 1072
rect 695 1038 707 1072
rect 583 1032 707 1038
rect 841 1072 965 1078
rect 841 1038 853 1072
rect 953 1038 965 1072
rect 841 1032 965 1038
rect 1099 1072 1223 1078
rect 1099 1038 1111 1072
rect 1211 1038 1223 1072
rect 1099 1032 1223 1038
rect 1357 1072 1481 1078
rect 1357 1038 1369 1072
rect 1469 1038 1481 1072
rect 1357 1032 1481 1038
rect 1615 1072 1739 1078
rect 1615 1038 1627 1072
rect 1727 1038 1739 1072
rect 1615 1032 1739 1038
rect 1873 1072 1997 1078
rect 1873 1038 1885 1072
rect 1985 1038 1997 1072
rect 1873 1032 1997 1038
rect 2131 1072 2255 1078
rect 2131 1038 2143 1072
rect 2243 1038 2255 1072
rect 2131 1032 2255 1038
rect 2389 1072 2513 1078
rect 2389 1038 2401 1072
rect 2501 1038 2513 1072
rect 2389 1032 2513 1038
rect 2647 1072 2771 1078
rect 2647 1038 2659 1072
rect 2759 1038 2771 1072
rect 2647 1032 2771 1038
rect 2905 1072 3029 1078
rect 2905 1038 2917 1072
rect 3017 1038 3029 1072
rect 2905 1032 3029 1038
rect 3163 1072 3287 1078
rect 3163 1038 3175 1072
rect 3275 1038 3287 1072
rect 3163 1032 3287 1038
rect 3421 1072 3545 1078
rect 3421 1038 3433 1072
rect 3533 1038 3545 1072
rect 3421 1032 3545 1038
rect 3679 1072 3803 1078
rect 3679 1038 3691 1072
rect 3791 1038 3803 1072
rect 3679 1032 3803 1038
rect 3937 1072 4061 1078
rect 3937 1038 3949 1072
rect 4049 1038 4061 1072
rect 3937 1032 4061 1038
rect 4195 1072 4319 1078
rect 4195 1038 4207 1072
rect 4307 1038 4319 1072
rect 4195 1032 4319 1038
rect -4409 988 -4363 1000
rect -4409 -988 -4403 988
rect -4369 -988 -4363 988
rect -4409 -1000 -4363 -988
rect -4151 988 -4105 1000
rect -4151 -988 -4145 988
rect -4111 -988 -4105 988
rect -4151 -1000 -4105 -988
rect -3893 988 -3847 1000
rect -3893 -988 -3887 988
rect -3853 -988 -3847 988
rect -3893 -1000 -3847 -988
rect -3635 988 -3589 1000
rect -3635 -988 -3629 988
rect -3595 -988 -3589 988
rect -3635 -1000 -3589 -988
rect -3377 988 -3331 1000
rect -3377 -988 -3371 988
rect -3337 -988 -3331 988
rect -3377 -1000 -3331 -988
rect -3119 988 -3073 1000
rect -3119 -988 -3113 988
rect -3079 -988 -3073 988
rect -3119 -1000 -3073 -988
rect -2861 988 -2815 1000
rect -2861 -988 -2855 988
rect -2821 -988 -2815 988
rect -2861 -1000 -2815 -988
rect -2603 988 -2557 1000
rect -2603 -988 -2597 988
rect -2563 -988 -2557 988
rect -2603 -1000 -2557 -988
rect -2345 988 -2299 1000
rect -2345 -988 -2339 988
rect -2305 -988 -2299 988
rect -2345 -1000 -2299 -988
rect -2087 988 -2041 1000
rect -2087 -988 -2081 988
rect -2047 -988 -2041 988
rect -2087 -1000 -2041 -988
rect -1829 988 -1783 1000
rect -1829 -988 -1823 988
rect -1789 -988 -1783 988
rect -1829 -1000 -1783 -988
rect -1571 988 -1525 1000
rect -1571 -988 -1565 988
rect -1531 -988 -1525 988
rect -1571 -1000 -1525 -988
rect -1313 988 -1267 1000
rect -1313 -988 -1307 988
rect -1273 -988 -1267 988
rect -1313 -1000 -1267 -988
rect -1055 988 -1009 1000
rect -1055 -988 -1049 988
rect -1015 -988 -1009 988
rect -1055 -1000 -1009 -988
rect -797 988 -751 1000
rect -797 -988 -791 988
rect -757 -988 -751 988
rect -797 -1000 -751 -988
rect -539 988 -493 1000
rect -539 -988 -533 988
rect -499 -988 -493 988
rect -539 -1000 -493 -988
rect -281 988 -235 1000
rect -281 -988 -275 988
rect -241 -988 -235 988
rect -281 -1000 -235 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 235 988 281 1000
rect 235 -988 241 988
rect 275 -988 281 988
rect 235 -1000 281 -988
rect 493 988 539 1000
rect 493 -988 499 988
rect 533 -988 539 988
rect 493 -1000 539 -988
rect 751 988 797 1000
rect 751 -988 757 988
rect 791 -988 797 988
rect 751 -1000 797 -988
rect 1009 988 1055 1000
rect 1009 -988 1015 988
rect 1049 -988 1055 988
rect 1009 -1000 1055 -988
rect 1267 988 1313 1000
rect 1267 -988 1273 988
rect 1307 -988 1313 988
rect 1267 -1000 1313 -988
rect 1525 988 1571 1000
rect 1525 -988 1531 988
rect 1565 -988 1571 988
rect 1525 -1000 1571 -988
rect 1783 988 1829 1000
rect 1783 -988 1789 988
rect 1823 -988 1829 988
rect 1783 -1000 1829 -988
rect 2041 988 2087 1000
rect 2041 -988 2047 988
rect 2081 -988 2087 988
rect 2041 -1000 2087 -988
rect 2299 988 2345 1000
rect 2299 -988 2305 988
rect 2339 -988 2345 988
rect 2299 -1000 2345 -988
rect 2557 988 2603 1000
rect 2557 -988 2563 988
rect 2597 -988 2603 988
rect 2557 -1000 2603 -988
rect 2815 988 2861 1000
rect 2815 -988 2821 988
rect 2855 -988 2861 988
rect 2815 -1000 2861 -988
rect 3073 988 3119 1000
rect 3073 -988 3079 988
rect 3113 -988 3119 988
rect 3073 -1000 3119 -988
rect 3331 988 3377 1000
rect 3331 -988 3337 988
rect 3371 -988 3377 988
rect 3331 -1000 3377 -988
rect 3589 988 3635 1000
rect 3589 -988 3595 988
rect 3629 -988 3635 988
rect 3589 -1000 3635 -988
rect 3847 988 3893 1000
rect 3847 -988 3853 988
rect 3887 -988 3893 988
rect 3847 -1000 3893 -988
rect 4105 988 4151 1000
rect 4105 -988 4111 988
rect 4145 -988 4151 988
rect 4105 -1000 4151 -988
rect 4363 988 4409 1000
rect 4363 -988 4369 988
rect 4403 -988 4409 988
rect 4363 -1000 4409 -988
rect -4319 -1038 -4195 -1032
rect -4319 -1072 -4307 -1038
rect -4207 -1072 -4195 -1038
rect -4319 -1078 -4195 -1072
rect -4061 -1038 -3937 -1032
rect -4061 -1072 -4049 -1038
rect -3949 -1072 -3937 -1038
rect -4061 -1078 -3937 -1072
rect -3803 -1038 -3679 -1032
rect -3803 -1072 -3791 -1038
rect -3691 -1072 -3679 -1038
rect -3803 -1078 -3679 -1072
rect -3545 -1038 -3421 -1032
rect -3545 -1072 -3533 -1038
rect -3433 -1072 -3421 -1038
rect -3545 -1078 -3421 -1072
rect -3287 -1038 -3163 -1032
rect -3287 -1072 -3275 -1038
rect -3175 -1072 -3163 -1038
rect -3287 -1078 -3163 -1072
rect -3029 -1038 -2905 -1032
rect -3029 -1072 -3017 -1038
rect -2917 -1072 -2905 -1038
rect -3029 -1078 -2905 -1072
rect -2771 -1038 -2647 -1032
rect -2771 -1072 -2759 -1038
rect -2659 -1072 -2647 -1038
rect -2771 -1078 -2647 -1072
rect -2513 -1038 -2389 -1032
rect -2513 -1072 -2501 -1038
rect -2401 -1072 -2389 -1038
rect -2513 -1078 -2389 -1072
rect -2255 -1038 -2131 -1032
rect -2255 -1072 -2243 -1038
rect -2143 -1072 -2131 -1038
rect -2255 -1078 -2131 -1072
rect -1997 -1038 -1873 -1032
rect -1997 -1072 -1985 -1038
rect -1885 -1072 -1873 -1038
rect -1997 -1078 -1873 -1072
rect -1739 -1038 -1615 -1032
rect -1739 -1072 -1727 -1038
rect -1627 -1072 -1615 -1038
rect -1739 -1078 -1615 -1072
rect -1481 -1038 -1357 -1032
rect -1481 -1072 -1469 -1038
rect -1369 -1072 -1357 -1038
rect -1481 -1078 -1357 -1072
rect -1223 -1038 -1099 -1032
rect -1223 -1072 -1211 -1038
rect -1111 -1072 -1099 -1038
rect -1223 -1078 -1099 -1072
rect -965 -1038 -841 -1032
rect -965 -1072 -953 -1038
rect -853 -1072 -841 -1038
rect -965 -1078 -841 -1072
rect -707 -1038 -583 -1032
rect -707 -1072 -695 -1038
rect -595 -1072 -583 -1038
rect -707 -1078 -583 -1072
rect -449 -1038 -325 -1032
rect -449 -1072 -437 -1038
rect -337 -1072 -325 -1038
rect -449 -1078 -325 -1072
rect -191 -1038 -67 -1032
rect -191 -1072 -179 -1038
rect -79 -1072 -67 -1038
rect -191 -1078 -67 -1072
rect 67 -1038 191 -1032
rect 67 -1072 79 -1038
rect 179 -1072 191 -1038
rect 67 -1078 191 -1072
rect 325 -1038 449 -1032
rect 325 -1072 337 -1038
rect 437 -1072 449 -1038
rect 325 -1078 449 -1072
rect 583 -1038 707 -1032
rect 583 -1072 595 -1038
rect 695 -1072 707 -1038
rect 583 -1078 707 -1072
rect 841 -1038 965 -1032
rect 841 -1072 853 -1038
rect 953 -1072 965 -1038
rect 841 -1078 965 -1072
rect 1099 -1038 1223 -1032
rect 1099 -1072 1111 -1038
rect 1211 -1072 1223 -1038
rect 1099 -1078 1223 -1072
rect 1357 -1038 1481 -1032
rect 1357 -1072 1369 -1038
rect 1469 -1072 1481 -1038
rect 1357 -1078 1481 -1072
rect 1615 -1038 1739 -1032
rect 1615 -1072 1627 -1038
rect 1727 -1072 1739 -1038
rect 1615 -1078 1739 -1072
rect 1873 -1038 1997 -1032
rect 1873 -1072 1885 -1038
rect 1985 -1072 1997 -1038
rect 1873 -1078 1997 -1072
rect 2131 -1038 2255 -1032
rect 2131 -1072 2143 -1038
rect 2243 -1072 2255 -1038
rect 2131 -1078 2255 -1072
rect 2389 -1038 2513 -1032
rect 2389 -1072 2401 -1038
rect 2501 -1072 2513 -1038
rect 2389 -1078 2513 -1072
rect 2647 -1038 2771 -1032
rect 2647 -1072 2659 -1038
rect 2759 -1072 2771 -1038
rect 2647 -1078 2771 -1072
rect 2905 -1038 3029 -1032
rect 2905 -1072 2917 -1038
rect 3017 -1072 3029 -1038
rect 2905 -1078 3029 -1072
rect 3163 -1038 3287 -1032
rect 3163 -1072 3175 -1038
rect 3275 -1072 3287 -1038
rect 3163 -1078 3287 -1072
rect 3421 -1038 3545 -1032
rect 3421 -1072 3433 -1038
rect 3533 -1072 3545 -1038
rect 3421 -1078 3545 -1072
rect 3679 -1038 3803 -1032
rect 3679 -1072 3691 -1038
rect 3791 -1072 3803 -1038
rect 3679 -1078 3803 -1072
rect 3937 -1038 4061 -1032
rect 3937 -1072 3949 -1038
rect 4049 -1072 4061 -1038
rect 3937 -1078 4061 -1072
rect 4195 -1038 4319 -1032
rect 4195 -1072 4207 -1038
rect 4307 -1072 4319 -1038
rect 4195 -1078 4319 -1072
<< properties >>
string FIXED_BBOX -4520 -1193 4520 1193
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10 l 1 m 1 nf 34 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713246000
<< pwell >>
rect -3405 -458 3405 458
<< mvnmos >>
rect -3177 -200 -2777 200
rect -2719 -200 -2319 200
rect -2261 -200 -1861 200
rect -1803 -200 -1403 200
rect -1345 -200 -945 200
rect -887 -200 -487 200
rect -429 -200 -29 200
rect 29 -200 429 200
rect 487 -200 887 200
rect 945 -200 1345 200
rect 1403 -200 1803 200
rect 1861 -200 2261 200
rect 2319 -200 2719 200
rect 2777 -200 3177 200
<< mvndiff >>
rect -3235 188 -3177 200
rect -3235 -188 -3223 188
rect -3189 -188 -3177 188
rect -3235 -200 -3177 -188
rect -2777 188 -2719 200
rect -2777 -188 -2765 188
rect -2731 -188 -2719 188
rect -2777 -200 -2719 -188
rect -2319 188 -2261 200
rect -2319 -188 -2307 188
rect -2273 -188 -2261 188
rect -2319 -200 -2261 -188
rect -1861 188 -1803 200
rect -1861 -188 -1849 188
rect -1815 -188 -1803 188
rect -1861 -200 -1803 -188
rect -1403 188 -1345 200
rect -1403 -188 -1391 188
rect -1357 -188 -1345 188
rect -1403 -200 -1345 -188
rect -945 188 -887 200
rect -945 -188 -933 188
rect -899 -188 -887 188
rect -945 -200 -887 -188
rect -487 188 -429 200
rect -487 -188 -475 188
rect -441 -188 -429 188
rect -487 -200 -429 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 429 188 487 200
rect 429 -188 441 188
rect 475 -188 487 188
rect 429 -200 487 -188
rect 887 188 945 200
rect 887 -188 899 188
rect 933 -188 945 188
rect 887 -200 945 -188
rect 1345 188 1403 200
rect 1345 -188 1357 188
rect 1391 -188 1403 188
rect 1345 -200 1403 -188
rect 1803 188 1861 200
rect 1803 -188 1815 188
rect 1849 -188 1861 188
rect 1803 -200 1861 -188
rect 2261 188 2319 200
rect 2261 -188 2273 188
rect 2307 -188 2319 188
rect 2261 -200 2319 -188
rect 2719 188 2777 200
rect 2719 -188 2731 188
rect 2765 -188 2777 188
rect 2719 -200 2777 -188
rect 3177 188 3235 200
rect 3177 -188 3189 188
rect 3223 -188 3235 188
rect 3177 -200 3235 -188
<< mvndiffc >>
rect -3223 -188 -3189 188
rect -2765 -188 -2731 188
rect -2307 -188 -2273 188
rect -1849 -188 -1815 188
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect 1815 -188 1849 188
rect 2273 -188 2307 188
rect 2731 -188 2765 188
rect 3189 -188 3223 188
<< mvpsubdiff >>
rect -3369 410 3369 422
rect -3369 376 -3261 410
rect 3261 376 3369 410
rect -3369 364 3369 376
rect -3369 314 -3311 364
rect -3369 -314 -3357 314
rect -3323 -314 -3311 314
rect 3311 314 3369 364
rect -3369 -364 -3311 -314
rect 3311 -314 3323 314
rect 3357 -314 3369 314
rect 3311 -364 3369 -314
rect -3369 -376 3369 -364
rect -3369 -410 -3261 -376
rect 3261 -410 3369 -376
rect -3369 -422 3369 -410
<< mvpsubdiffcont >>
rect -3261 376 3261 410
rect -3357 -314 -3323 314
rect 3323 -314 3357 314
rect -3261 -410 3261 -376
<< poly >>
rect -3122 272 -2832 288
rect -3122 255 -3106 272
rect -3177 238 -3106 255
rect -2848 255 -2832 272
rect -2664 272 -2374 288
rect -2664 255 -2648 272
rect -2848 238 -2777 255
rect -3177 200 -2777 238
rect -2719 238 -2648 255
rect -2390 255 -2374 272
rect -2206 272 -1916 288
rect -2206 255 -2190 272
rect -2390 238 -2319 255
rect -2719 200 -2319 238
rect -2261 238 -2190 255
rect -1932 255 -1916 272
rect -1748 272 -1458 288
rect -1748 255 -1732 272
rect -1932 238 -1861 255
rect -2261 200 -1861 238
rect -1803 238 -1732 255
rect -1474 255 -1458 272
rect -1290 272 -1000 288
rect -1290 255 -1274 272
rect -1474 238 -1403 255
rect -1803 200 -1403 238
rect -1345 238 -1274 255
rect -1016 255 -1000 272
rect -832 272 -542 288
rect -832 255 -816 272
rect -1016 238 -945 255
rect -1345 200 -945 238
rect -887 238 -816 255
rect -558 255 -542 272
rect -374 272 -84 288
rect -374 255 -358 272
rect -558 238 -487 255
rect -887 200 -487 238
rect -429 238 -358 255
rect -100 255 -84 272
rect 84 272 374 288
rect 84 255 100 272
rect -100 238 -29 255
rect -429 200 -29 238
rect 29 238 100 255
rect 358 255 374 272
rect 542 272 832 288
rect 542 255 558 272
rect 358 238 429 255
rect 29 200 429 238
rect 487 238 558 255
rect 816 255 832 272
rect 1000 272 1290 288
rect 1000 255 1016 272
rect 816 238 887 255
rect 487 200 887 238
rect 945 238 1016 255
rect 1274 255 1290 272
rect 1458 272 1748 288
rect 1458 255 1474 272
rect 1274 238 1345 255
rect 945 200 1345 238
rect 1403 238 1474 255
rect 1732 255 1748 272
rect 1916 272 2206 288
rect 1916 255 1932 272
rect 1732 238 1803 255
rect 1403 200 1803 238
rect 1861 238 1932 255
rect 2190 255 2206 272
rect 2374 272 2664 288
rect 2374 255 2390 272
rect 2190 238 2261 255
rect 1861 200 2261 238
rect 2319 238 2390 255
rect 2648 255 2664 272
rect 2832 272 3122 288
rect 2832 255 2848 272
rect 2648 238 2719 255
rect 2319 200 2719 238
rect 2777 238 2848 255
rect 3106 255 3122 272
rect 3106 238 3177 255
rect 2777 200 3177 238
rect -3177 -238 -2777 -200
rect -3177 -255 -3106 -238
rect -3122 -272 -3106 -255
rect -2848 -255 -2777 -238
rect -2719 -238 -2319 -200
rect -2719 -255 -2648 -238
rect -2848 -272 -2832 -255
rect -3122 -288 -2832 -272
rect -2664 -272 -2648 -255
rect -2390 -255 -2319 -238
rect -2261 -238 -1861 -200
rect -2261 -255 -2190 -238
rect -2390 -272 -2374 -255
rect -2664 -288 -2374 -272
rect -2206 -272 -2190 -255
rect -1932 -255 -1861 -238
rect -1803 -238 -1403 -200
rect -1803 -255 -1732 -238
rect -1932 -272 -1916 -255
rect -2206 -288 -1916 -272
rect -1748 -272 -1732 -255
rect -1474 -255 -1403 -238
rect -1345 -238 -945 -200
rect -1345 -255 -1274 -238
rect -1474 -272 -1458 -255
rect -1748 -288 -1458 -272
rect -1290 -272 -1274 -255
rect -1016 -255 -945 -238
rect -887 -238 -487 -200
rect -887 -255 -816 -238
rect -1016 -272 -1000 -255
rect -1290 -288 -1000 -272
rect -832 -272 -816 -255
rect -558 -255 -487 -238
rect -429 -238 -29 -200
rect -429 -255 -358 -238
rect -558 -272 -542 -255
rect -832 -288 -542 -272
rect -374 -272 -358 -255
rect -100 -255 -29 -238
rect 29 -238 429 -200
rect 29 -255 100 -238
rect -100 -272 -84 -255
rect -374 -288 -84 -272
rect 84 -272 100 -255
rect 358 -255 429 -238
rect 487 -238 887 -200
rect 487 -255 558 -238
rect 358 -272 374 -255
rect 84 -288 374 -272
rect 542 -272 558 -255
rect 816 -255 887 -238
rect 945 -238 1345 -200
rect 945 -255 1016 -238
rect 816 -272 832 -255
rect 542 -288 832 -272
rect 1000 -272 1016 -255
rect 1274 -255 1345 -238
rect 1403 -238 1803 -200
rect 1403 -255 1474 -238
rect 1274 -272 1290 -255
rect 1000 -288 1290 -272
rect 1458 -272 1474 -255
rect 1732 -255 1803 -238
rect 1861 -238 2261 -200
rect 1861 -255 1932 -238
rect 1732 -272 1748 -255
rect 1458 -288 1748 -272
rect 1916 -272 1932 -255
rect 2190 -255 2261 -238
rect 2319 -238 2719 -200
rect 2319 -255 2390 -238
rect 2190 -272 2206 -255
rect 1916 -288 2206 -272
rect 2374 -272 2390 -255
rect 2648 -255 2719 -238
rect 2777 -238 3177 -200
rect 2777 -255 2848 -238
rect 2648 -272 2664 -255
rect 2374 -288 2664 -272
rect 2832 -272 2848 -255
rect 3106 -255 3177 -238
rect 3106 -272 3122 -255
rect 2832 -288 3122 -272
<< polycont >>
rect -3106 238 -2848 272
rect -2648 238 -2390 272
rect -2190 238 -1932 272
rect -1732 238 -1474 272
rect -1274 238 -1016 272
rect -816 238 -558 272
rect -358 238 -100 272
rect 100 238 358 272
rect 558 238 816 272
rect 1016 238 1274 272
rect 1474 238 1732 272
rect 1932 238 2190 272
rect 2390 238 2648 272
rect 2848 238 3106 272
rect -3106 -272 -2848 -238
rect -2648 -272 -2390 -238
rect -2190 -272 -1932 -238
rect -1732 -272 -1474 -238
rect -1274 -272 -1016 -238
rect -816 -272 -558 -238
rect -358 -272 -100 -238
rect 100 -272 358 -238
rect 558 -272 816 -238
rect 1016 -272 1274 -238
rect 1474 -272 1732 -238
rect 1932 -272 2190 -238
rect 2390 -272 2648 -238
rect 2848 -272 3106 -238
<< locali >>
rect -3357 376 -3261 410
rect 3261 376 3357 410
rect -3357 314 -3323 376
rect 3323 314 3357 376
rect -3122 238 -3106 272
rect -2848 238 -2832 272
rect -2664 238 -2648 272
rect -2390 238 -2374 272
rect -2206 238 -2190 272
rect -1932 238 -1916 272
rect -1748 238 -1732 272
rect -1474 238 -1458 272
rect -1290 238 -1274 272
rect -1016 238 -1000 272
rect -832 238 -816 272
rect -558 238 -542 272
rect -374 238 -358 272
rect -100 238 -84 272
rect 84 238 100 272
rect 358 238 374 272
rect 542 238 558 272
rect 816 238 832 272
rect 1000 238 1016 272
rect 1274 238 1290 272
rect 1458 238 1474 272
rect 1732 238 1748 272
rect 1916 238 1932 272
rect 2190 238 2206 272
rect 2374 238 2390 272
rect 2648 238 2664 272
rect 2832 238 2848 272
rect 3106 238 3122 272
rect -3223 188 -3189 204
rect -3223 -204 -3189 -188
rect -2765 188 -2731 204
rect -2765 -204 -2731 -188
rect -2307 188 -2273 204
rect -2307 -204 -2273 -188
rect -1849 188 -1815 204
rect -1849 -204 -1815 -188
rect -1391 188 -1357 204
rect -1391 -204 -1357 -188
rect -933 188 -899 204
rect -933 -204 -899 -188
rect -475 188 -441 204
rect -475 -204 -441 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 441 188 475 204
rect 441 -204 475 -188
rect 899 188 933 204
rect 899 -204 933 -188
rect 1357 188 1391 204
rect 1357 -204 1391 -188
rect 1815 188 1849 204
rect 1815 -204 1849 -188
rect 2273 188 2307 204
rect 2273 -204 2307 -188
rect 2731 188 2765 204
rect 2731 -204 2765 -188
rect 3189 188 3223 204
rect 3189 -204 3223 -188
rect -3122 -272 -3106 -238
rect -2848 -272 -2832 -238
rect -2664 -272 -2648 -238
rect -2390 -272 -2374 -238
rect -2206 -272 -2190 -238
rect -1932 -272 -1916 -238
rect -1748 -272 -1732 -238
rect -1474 -272 -1458 -238
rect -1290 -272 -1274 -238
rect -1016 -272 -1000 -238
rect -832 -272 -816 -238
rect -558 -272 -542 -238
rect -374 -272 -358 -238
rect -100 -272 -84 -238
rect 84 -272 100 -238
rect 358 -272 374 -238
rect 542 -272 558 -238
rect 816 -272 832 -238
rect 1000 -272 1016 -238
rect 1274 -272 1290 -238
rect 1458 -272 1474 -238
rect 1732 -272 1748 -238
rect 1916 -272 1932 -238
rect 2190 -272 2206 -238
rect 2374 -272 2390 -238
rect 2648 -272 2664 -238
rect 2832 -272 2848 -238
rect 3106 -272 3122 -238
rect -3357 -376 -3323 -314
rect 3323 -376 3357 -314
rect -3357 -410 -3261 -376
rect 3261 -410 3357 -376
<< viali >>
rect -3106 238 -2848 272
rect -2648 238 -2390 272
rect -2190 238 -1932 272
rect -1732 238 -1474 272
rect -1274 238 -1016 272
rect -816 238 -558 272
rect -358 238 -100 272
rect 100 238 358 272
rect 558 238 816 272
rect 1016 238 1274 272
rect 1474 238 1732 272
rect 1932 238 2190 272
rect 2390 238 2648 272
rect 2848 238 3106 272
rect -3223 -188 -3189 188
rect -2765 -188 -2731 188
rect -2307 -188 -2273 188
rect -1849 -188 -1815 188
rect -1391 -188 -1357 188
rect -933 -188 -899 188
rect -475 -188 -441 188
rect -17 -188 17 188
rect 441 -188 475 188
rect 899 -188 933 188
rect 1357 -188 1391 188
rect 1815 -188 1849 188
rect 2273 -188 2307 188
rect 2731 -188 2765 188
rect 3189 -188 3223 188
rect -3106 -272 -2848 -238
rect -2648 -272 -2390 -238
rect -2190 -272 -1932 -238
rect -1732 -272 -1474 -238
rect -1274 -272 -1016 -238
rect -816 -272 -558 -238
rect -358 -272 -100 -238
rect 100 -272 358 -238
rect 558 -272 816 -238
rect 1016 -272 1274 -238
rect 1474 -272 1732 -238
rect 1932 -272 2190 -238
rect 2390 -272 2648 -238
rect 2848 -272 3106 -238
<< metal1 >>
rect -3118 272 -2836 278
rect -3118 238 -3106 272
rect -2848 238 -2836 272
rect -3118 232 -2836 238
rect -2660 272 -2378 278
rect -2660 238 -2648 272
rect -2390 238 -2378 272
rect -2660 232 -2378 238
rect -2202 272 -1920 278
rect -2202 238 -2190 272
rect -1932 238 -1920 272
rect -2202 232 -1920 238
rect -1744 272 -1462 278
rect -1744 238 -1732 272
rect -1474 238 -1462 272
rect -1744 232 -1462 238
rect -1286 272 -1004 278
rect -1286 238 -1274 272
rect -1016 238 -1004 272
rect -1286 232 -1004 238
rect -828 272 -546 278
rect -828 238 -816 272
rect -558 238 -546 272
rect -828 232 -546 238
rect -370 272 -88 278
rect -370 238 -358 272
rect -100 238 -88 272
rect -370 232 -88 238
rect 88 272 370 278
rect 88 238 100 272
rect 358 238 370 272
rect 88 232 370 238
rect 546 272 828 278
rect 546 238 558 272
rect 816 238 828 272
rect 546 232 828 238
rect 1004 272 1286 278
rect 1004 238 1016 272
rect 1274 238 1286 272
rect 1004 232 1286 238
rect 1462 272 1744 278
rect 1462 238 1474 272
rect 1732 238 1744 272
rect 1462 232 1744 238
rect 1920 272 2202 278
rect 1920 238 1932 272
rect 2190 238 2202 272
rect 1920 232 2202 238
rect 2378 272 2660 278
rect 2378 238 2390 272
rect 2648 238 2660 272
rect 2378 232 2660 238
rect 2836 272 3118 278
rect 2836 238 2848 272
rect 3106 238 3118 272
rect 2836 232 3118 238
rect -3229 188 -3183 200
rect -3229 -188 -3223 188
rect -3189 -188 -3183 188
rect -3229 -200 -3183 -188
rect -2771 188 -2725 200
rect -2771 -188 -2765 188
rect -2731 -188 -2725 188
rect -2771 -200 -2725 -188
rect -2313 188 -2267 200
rect -2313 -188 -2307 188
rect -2273 -188 -2267 188
rect -2313 -200 -2267 -188
rect -1855 188 -1809 200
rect -1855 -188 -1849 188
rect -1815 -188 -1809 188
rect -1855 -200 -1809 -188
rect -1397 188 -1351 200
rect -1397 -188 -1391 188
rect -1357 -188 -1351 188
rect -1397 -200 -1351 -188
rect -939 188 -893 200
rect -939 -188 -933 188
rect -899 -188 -893 188
rect -939 -200 -893 -188
rect -481 188 -435 200
rect -481 -188 -475 188
rect -441 -188 -435 188
rect -481 -200 -435 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 435 188 481 200
rect 435 -188 441 188
rect 475 -188 481 188
rect 435 -200 481 -188
rect 893 188 939 200
rect 893 -188 899 188
rect 933 -188 939 188
rect 893 -200 939 -188
rect 1351 188 1397 200
rect 1351 -188 1357 188
rect 1391 -188 1397 188
rect 1351 -200 1397 -188
rect 1809 188 1855 200
rect 1809 -188 1815 188
rect 1849 -188 1855 188
rect 1809 -200 1855 -188
rect 2267 188 2313 200
rect 2267 -188 2273 188
rect 2307 -188 2313 188
rect 2267 -200 2313 -188
rect 2725 188 2771 200
rect 2725 -188 2731 188
rect 2765 -188 2771 188
rect 2725 -200 2771 -188
rect 3183 188 3229 200
rect 3183 -188 3189 188
rect 3223 -188 3229 188
rect 3183 -200 3229 -188
rect -3118 -238 -2836 -232
rect -3118 -272 -3106 -238
rect -2848 -272 -2836 -238
rect -3118 -278 -2836 -272
rect -2660 -238 -2378 -232
rect -2660 -272 -2648 -238
rect -2390 -272 -2378 -238
rect -2660 -278 -2378 -272
rect -2202 -238 -1920 -232
rect -2202 -272 -2190 -238
rect -1932 -272 -1920 -238
rect -2202 -278 -1920 -272
rect -1744 -238 -1462 -232
rect -1744 -272 -1732 -238
rect -1474 -272 -1462 -238
rect -1744 -278 -1462 -272
rect -1286 -238 -1004 -232
rect -1286 -272 -1274 -238
rect -1016 -272 -1004 -238
rect -1286 -278 -1004 -272
rect -828 -238 -546 -232
rect -828 -272 -816 -238
rect -558 -272 -546 -238
rect -828 -278 -546 -272
rect -370 -238 -88 -232
rect -370 -272 -358 -238
rect -100 -272 -88 -238
rect -370 -278 -88 -272
rect 88 -238 370 -232
rect 88 -272 100 -238
rect 358 -272 370 -238
rect 88 -278 370 -272
rect 546 -238 828 -232
rect 546 -272 558 -238
rect 816 -272 828 -238
rect 546 -278 828 -272
rect 1004 -238 1286 -232
rect 1004 -272 1016 -238
rect 1274 -272 1286 -238
rect 1004 -278 1286 -272
rect 1462 -238 1744 -232
rect 1462 -272 1474 -238
rect 1732 -272 1744 -238
rect 1462 -278 1744 -272
rect 1920 -238 2202 -232
rect 1920 -272 1932 -238
rect 2190 -272 2202 -238
rect 1920 -278 2202 -272
rect 2378 -238 2660 -232
rect 2378 -272 2390 -238
rect 2648 -272 2660 -238
rect 2378 -278 2660 -272
rect 2836 -238 3118 -232
rect 2836 -272 2848 -238
rect 3106 -272 3118 -238
rect 2836 -278 3118 -272
<< properties >>
string FIXED_BBOX -3340 -393 3340 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 2 m 1 nf 14 diffcov 100 polycov 70 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

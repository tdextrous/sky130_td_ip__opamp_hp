magic
tech sky130A
magscale 1 2
timestamp 1713285936
<< pwell >>
rect -5359 -458 5359 458
<< mvnmos >>
rect -5131 -200 -4931 200
rect -4873 -200 -4673 200
rect -4615 -200 -4415 200
rect -4357 -200 -4157 200
rect -4099 -200 -3899 200
rect -3841 -200 -3641 200
rect -3583 -200 -3383 200
rect -3325 -200 -3125 200
rect -3067 -200 -2867 200
rect -2809 -200 -2609 200
rect -2551 -200 -2351 200
rect -2293 -200 -2093 200
rect -2035 -200 -1835 200
rect -1777 -200 -1577 200
rect -1519 -200 -1319 200
rect -1261 -200 -1061 200
rect -1003 -200 -803 200
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
rect 803 -200 1003 200
rect 1061 -200 1261 200
rect 1319 -200 1519 200
rect 1577 -200 1777 200
rect 1835 -200 2035 200
rect 2093 -200 2293 200
rect 2351 -200 2551 200
rect 2609 -200 2809 200
rect 2867 -200 3067 200
rect 3125 -200 3325 200
rect 3383 -200 3583 200
rect 3641 -200 3841 200
rect 3899 -200 4099 200
rect 4157 -200 4357 200
rect 4415 -200 4615 200
rect 4673 -200 4873 200
rect 4931 -200 5131 200
<< mvndiff >>
rect -5189 188 -5131 200
rect -5189 -188 -5177 188
rect -5143 -188 -5131 188
rect -5189 -200 -5131 -188
rect -4931 188 -4873 200
rect -4931 -188 -4919 188
rect -4885 -188 -4873 188
rect -4931 -200 -4873 -188
rect -4673 188 -4615 200
rect -4673 -188 -4661 188
rect -4627 -188 -4615 188
rect -4673 -200 -4615 -188
rect -4415 188 -4357 200
rect -4415 -188 -4403 188
rect -4369 -188 -4357 188
rect -4415 -200 -4357 -188
rect -4157 188 -4099 200
rect -4157 -188 -4145 188
rect -4111 -188 -4099 188
rect -4157 -200 -4099 -188
rect -3899 188 -3841 200
rect -3899 -188 -3887 188
rect -3853 -188 -3841 188
rect -3899 -200 -3841 -188
rect -3641 188 -3583 200
rect -3641 -188 -3629 188
rect -3595 -188 -3583 188
rect -3641 -200 -3583 -188
rect -3383 188 -3325 200
rect -3383 -188 -3371 188
rect -3337 -188 -3325 188
rect -3383 -200 -3325 -188
rect -3125 188 -3067 200
rect -3125 -188 -3113 188
rect -3079 -188 -3067 188
rect -3125 -200 -3067 -188
rect -2867 188 -2809 200
rect -2867 -188 -2855 188
rect -2821 -188 -2809 188
rect -2867 -200 -2809 -188
rect -2609 188 -2551 200
rect -2609 -188 -2597 188
rect -2563 -188 -2551 188
rect -2609 -200 -2551 -188
rect -2351 188 -2293 200
rect -2351 -188 -2339 188
rect -2305 -188 -2293 188
rect -2351 -200 -2293 -188
rect -2093 188 -2035 200
rect -2093 -188 -2081 188
rect -2047 -188 -2035 188
rect -2093 -200 -2035 -188
rect -1835 188 -1777 200
rect -1835 -188 -1823 188
rect -1789 -188 -1777 188
rect -1835 -200 -1777 -188
rect -1577 188 -1519 200
rect -1577 -188 -1565 188
rect -1531 -188 -1519 188
rect -1577 -200 -1519 -188
rect -1319 188 -1261 200
rect -1319 -188 -1307 188
rect -1273 -188 -1261 188
rect -1319 -200 -1261 -188
rect -1061 188 -1003 200
rect -1061 -188 -1049 188
rect -1015 -188 -1003 188
rect -1061 -200 -1003 -188
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
rect 1003 188 1061 200
rect 1003 -188 1015 188
rect 1049 -188 1061 188
rect 1003 -200 1061 -188
rect 1261 188 1319 200
rect 1261 -188 1273 188
rect 1307 -188 1319 188
rect 1261 -200 1319 -188
rect 1519 188 1577 200
rect 1519 -188 1531 188
rect 1565 -188 1577 188
rect 1519 -200 1577 -188
rect 1777 188 1835 200
rect 1777 -188 1789 188
rect 1823 -188 1835 188
rect 1777 -200 1835 -188
rect 2035 188 2093 200
rect 2035 -188 2047 188
rect 2081 -188 2093 188
rect 2035 -200 2093 -188
rect 2293 188 2351 200
rect 2293 -188 2305 188
rect 2339 -188 2351 188
rect 2293 -200 2351 -188
rect 2551 188 2609 200
rect 2551 -188 2563 188
rect 2597 -188 2609 188
rect 2551 -200 2609 -188
rect 2809 188 2867 200
rect 2809 -188 2821 188
rect 2855 -188 2867 188
rect 2809 -200 2867 -188
rect 3067 188 3125 200
rect 3067 -188 3079 188
rect 3113 -188 3125 188
rect 3067 -200 3125 -188
rect 3325 188 3383 200
rect 3325 -188 3337 188
rect 3371 -188 3383 188
rect 3325 -200 3383 -188
rect 3583 188 3641 200
rect 3583 -188 3595 188
rect 3629 -188 3641 188
rect 3583 -200 3641 -188
rect 3841 188 3899 200
rect 3841 -188 3853 188
rect 3887 -188 3899 188
rect 3841 -200 3899 -188
rect 4099 188 4157 200
rect 4099 -188 4111 188
rect 4145 -188 4157 188
rect 4099 -200 4157 -188
rect 4357 188 4415 200
rect 4357 -188 4369 188
rect 4403 -188 4415 188
rect 4357 -200 4415 -188
rect 4615 188 4673 200
rect 4615 -188 4627 188
rect 4661 -188 4673 188
rect 4615 -200 4673 -188
rect 4873 188 4931 200
rect 4873 -188 4885 188
rect 4919 -188 4931 188
rect 4873 -200 4931 -188
rect 5131 188 5189 200
rect 5131 -188 5143 188
rect 5177 -188 5189 188
rect 5131 -200 5189 -188
<< mvndiffc >>
rect -5177 -188 -5143 188
rect -4919 -188 -4885 188
rect -4661 -188 -4627 188
rect -4403 -188 -4369 188
rect -4145 -188 -4111 188
rect -3887 -188 -3853 188
rect -3629 -188 -3595 188
rect -3371 -188 -3337 188
rect -3113 -188 -3079 188
rect -2855 -188 -2821 188
rect -2597 -188 -2563 188
rect -2339 -188 -2305 188
rect -2081 -188 -2047 188
rect -1823 -188 -1789 188
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect 1789 -188 1823 188
rect 2047 -188 2081 188
rect 2305 -188 2339 188
rect 2563 -188 2597 188
rect 2821 -188 2855 188
rect 3079 -188 3113 188
rect 3337 -188 3371 188
rect 3595 -188 3629 188
rect 3853 -188 3887 188
rect 4111 -188 4145 188
rect 4369 -188 4403 188
rect 4627 -188 4661 188
rect 4885 -188 4919 188
rect 5143 -188 5177 188
<< mvpsubdiff >>
rect -5323 410 5323 422
rect -5323 376 -5215 410
rect 5215 376 5323 410
rect -5323 364 5323 376
rect -5323 314 -5265 364
rect -5323 -314 -5311 314
rect -5277 -314 -5265 314
rect 5265 314 5323 364
rect -5323 -364 -5265 -314
rect 5265 -314 5277 314
rect 5311 -314 5323 314
rect 5265 -364 5323 -314
rect -5323 -376 5323 -364
rect -5323 -410 -5215 -376
rect 5215 -410 5323 -376
rect -5323 -422 5323 -410
<< mvpsubdiffcont >>
rect -5215 376 5215 410
rect -5311 -314 -5277 314
rect 5277 -314 5311 314
rect -5215 -410 5215 -376
<< poly >>
rect -5097 272 -4965 288
rect -5097 255 -5081 272
rect -5131 238 -5081 255
rect -4981 255 -4965 272
rect -4839 272 -4707 288
rect -4839 255 -4823 272
rect -4981 238 -4931 255
rect -5131 200 -4931 238
rect -4873 238 -4823 255
rect -4723 255 -4707 272
rect -4581 272 -4449 288
rect -4581 255 -4565 272
rect -4723 238 -4673 255
rect -4873 200 -4673 238
rect -4615 238 -4565 255
rect -4465 255 -4449 272
rect -4323 272 -4191 288
rect -4323 255 -4307 272
rect -4465 238 -4415 255
rect -4615 200 -4415 238
rect -4357 238 -4307 255
rect -4207 255 -4191 272
rect -4065 272 -3933 288
rect -4065 255 -4049 272
rect -4207 238 -4157 255
rect -4357 200 -4157 238
rect -4099 238 -4049 255
rect -3949 255 -3933 272
rect -3807 272 -3675 288
rect -3807 255 -3791 272
rect -3949 238 -3899 255
rect -4099 200 -3899 238
rect -3841 238 -3791 255
rect -3691 255 -3675 272
rect -3549 272 -3417 288
rect -3549 255 -3533 272
rect -3691 238 -3641 255
rect -3841 200 -3641 238
rect -3583 238 -3533 255
rect -3433 255 -3417 272
rect -3291 272 -3159 288
rect -3291 255 -3275 272
rect -3433 238 -3383 255
rect -3583 200 -3383 238
rect -3325 238 -3275 255
rect -3175 255 -3159 272
rect -3033 272 -2901 288
rect -3033 255 -3017 272
rect -3175 238 -3125 255
rect -3325 200 -3125 238
rect -3067 238 -3017 255
rect -2917 255 -2901 272
rect -2775 272 -2643 288
rect -2775 255 -2759 272
rect -2917 238 -2867 255
rect -3067 200 -2867 238
rect -2809 238 -2759 255
rect -2659 255 -2643 272
rect -2517 272 -2385 288
rect -2517 255 -2501 272
rect -2659 238 -2609 255
rect -2809 200 -2609 238
rect -2551 238 -2501 255
rect -2401 255 -2385 272
rect -2259 272 -2127 288
rect -2259 255 -2243 272
rect -2401 238 -2351 255
rect -2551 200 -2351 238
rect -2293 238 -2243 255
rect -2143 255 -2127 272
rect -2001 272 -1869 288
rect -2001 255 -1985 272
rect -2143 238 -2093 255
rect -2293 200 -2093 238
rect -2035 238 -1985 255
rect -1885 255 -1869 272
rect -1743 272 -1611 288
rect -1743 255 -1727 272
rect -1885 238 -1835 255
rect -2035 200 -1835 238
rect -1777 238 -1727 255
rect -1627 255 -1611 272
rect -1485 272 -1353 288
rect -1485 255 -1469 272
rect -1627 238 -1577 255
rect -1777 200 -1577 238
rect -1519 238 -1469 255
rect -1369 255 -1353 272
rect -1227 272 -1095 288
rect -1227 255 -1211 272
rect -1369 238 -1319 255
rect -1519 200 -1319 238
rect -1261 238 -1211 255
rect -1111 255 -1095 272
rect -969 272 -837 288
rect -969 255 -953 272
rect -1111 238 -1061 255
rect -1261 200 -1061 238
rect -1003 238 -953 255
rect -853 255 -837 272
rect -711 272 -579 288
rect -711 255 -695 272
rect -853 238 -803 255
rect -1003 200 -803 238
rect -745 238 -695 255
rect -595 255 -579 272
rect -453 272 -321 288
rect -453 255 -437 272
rect -595 238 -545 255
rect -745 200 -545 238
rect -487 238 -437 255
rect -337 255 -321 272
rect -195 272 -63 288
rect -195 255 -179 272
rect -337 238 -287 255
rect -487 200 -287 238
rect -229 238 -179 255
rect -79 255 -63 272
rect 63 272 195 288
rect 63 255 79 272
rect -79 238 -29 255
rect -229 200 -29 238
rect 29 238 79 255
rect 179 255 195 272
rect 321 272 453 288
rect 321 255 337 272
rect 179 238 229 255
rect 29 200 229 238
rect 287 238 337 255
rect 437 255 453 272
rect 579 272 711 288
rect 579 255 595 272
rect 437 238 487 255
rect 287 200 487 238
rect 545 238 595 255
rect 695 255 711 272
rect 837 272 969 288
rect 837 255 853 272
rect 695 238 745 255
rect 545 200 745 238
rect 803 238 853 255
rect 953 255 969 272
rect 1095 272 1227 288
rect 1095 255 1111 272
rect 953 238 1003 255
rect 803 200 1003 238
rect 1061 238 1111 255
rect 1211 255 1227 272
rect 1353 272 1485 288
rect 1353 255 1369 272
rect 1211 238 1261 255
rect 1061 200 1261 238
rect 1319 238 1369 255
rect 1469 255 1485 272
rect 1611 272 1743 288
rect 1611 255 1627 272
rect 1469 238 1519 255
rect 1319 200 1519 238
rect 1577 238 1627 255
rect 1727 255 1743 272
rect 1869 272 2001 288
rect 1869 255 1885 272
rect 1727 238 1777 255
rect 1577 200 1777 238
rect 1835 238 1885 255
rect 1985 255 2001 272
rect 2127 272 2259 288
rect 2127 255 2143 272
rect 1985 238 2035 255
rect 1835 200 2035 238
rect 2093 238 2143 255
rect 2243 255 2259 272
rect 2385 272 2517 288
rect 2385 255 2401 272
rect 2243 238 2293 255
rect 2093 200 2293 238
rect 2351 238 2401 255
rect 2501 255 2517 272
rect 2643 272 2775 288
rect 2643 255 2659 272
rect 2501 238 2551 255
rect 2351 200 2551 238
rect 2609 238 2659 255
rect 2759 255 2775 272
rect 2901 272 3033 288
rect 2901 255 2917 272
rect 2759 238 2809 255
rect 2609 200 2809 238
rect 2867 238 2917 255
rect 3017 255 3033 272
rect 3159 272 3291 288
rect 3159 255 3175 272
rect 3017 238 3067 255
rect 2867 200 3067 238
rect 3125 238 3175 255
rect 3275 255 3291 272
rect 3417 272 3549 288
rect 3417 255 3433 272
rect 3275 238 3325 255
rect 3125 200 3325 238
rect 3383 238 3433 255
rect 3533 255 3549 272
rect 3675 272 3807 288
rect 3675 255 3691 272
rect 3533 238 3583 255
rect 3383 200 3583 238
rect 3641 238 3691 255
rect 3791 255 3807 272
rect 3933 272 4065 288
rect 3933 255 3949 272
rect 3791 238 3841 255
rect 3641 200 3841 238
rect 3899 238 3949 255
rect 4049 255 4065 272
rect 4191 272 4323 288
rect 4191 255 4207 272
rect 4049 238 4099 255
rect 3899 200 4099 238
rect 4157 238 4207 255
rect 4307 255 4323 272
rect 4449 272 4581 288
rect 4449 255 4465 272
rect 4307 238 4357 255
rect 4157 200 4357 238
rect 4415 238 4465 255
rect 4565 255 4581 272
rect 4707 272 4839 288
rect 4707 255 4723 272
rect 4565 238 4615 255
rect 4415 200 4615 238
rect 4673 238 4723 255
rect 4823 255 4839 272
rect 4965 272 5097 288
rect 4965 255 4981 272
rect 4823 238 4873 255
rect 4673 200 4873 238
rect 4931 238 4981 255
rect 5081 255 5097 272
rect 5081 238 5131 255
rect 4931 200 5131 238
rect -5131 -238 -4931 -200
rect -5131 -255 -5081 -238
rect -5097 -272 -5081 -255
rect -4981 -255 -4931 -238
rect -4873 -238 -4673 -200
rect -4873 -255 -4823 -238
rect -4981 -272 -4965 -255
rect -5097 -288 -4965 -272
rect -4839 -272 -4823 -255
rect -4723 -255 -4673 -238
rect -4615 -238 -4415 -200
rect -4615 -255 -4565 -238
rect -4723 -272 -4707 -255
rect -4839 -288 -4707 -272
rect -4581 -272 -4565 -255
rect -4465 -255 -4415 -238
rect -4357 -238 -4157 -200
rect -4357 -255 -4307 -238
rect -4465 -272 -4449 -255
rect -4581 -288 -4449 -272
rect -4323 -272 -4307 -255
rect -4207 -255 -4157 -238
rect -4099 -238 -3899 -200
rect -4099 -255 -4049 -238
rect -4207 -272 -4191 -255
rect -4323 -288 -4191 -272
rect -4065 -272 -4049 -255
rect -3949 -255 -3899 -238
rect -3841 -238 -3641 -200
rect -3841 -255 -3791 -238
rect -3949 -272 -3933 -255
rect -4065 -288 -3933 -272
rect -3807 -272 -3791 -255
rect -3691 -255 -3641 -238
rect -3583 -238 -3383 -200
rect -3583 -255 -3533 -238
rect -3691 -272 -3675 -255
rect -3807 -288 -3675 -272
rect -3549 -272 -3533 -255
rect -3433 -255 -3383 -238
rect -3325 -238 -3125 -200
rect -3325 -255 -3275 -238
rect -3433 -272 -3417 -255
rect -3549 -288 -3417 -272
rect -3291 -272 -3275 -255
rect -3175 -255 -3125 -238
rect -3067 -238 -2867 -200
rect -3067 -255 -3017 -238
rect -3175 -272 -3159 -255
rect -3291 -288 -3159 -272
rect -3033 -272 -3017 -255
rect -2917 -255 -2867 -238
rect -2809 -238 -2609 -200
rect -2809 -255 -2759 -238
rect -2917 -272 -2901 -255
rect -3033 -288 -2901 -272
rect -2775 -272 -2759 -255
rect -2659 -255 -2609 -238
rect -2551 -238 -2351 -200
rect -2551 -255 -2501 -238
rect -2659 -272 -2643 -255
rect -2775 -288 -2643 -272
rect -2517 -272 -2501 -255
rect -2401 -255 -2351 -238
rect -2293 -238 -2093 -200
rect -2293 -255 -2243 -238
rect -2401 -272 -2385 -255
rect -2517 -288 -2385 -272
rect -2259 -272 -2243 -255
rect -2143 -255 -2093 -238
rect -2035 -238 -1835 -200
rect -2035 -255 -1985 -238
rect -2143 -272 -2127 -255
rect -2259 -288 -2127 -272
rect -2001 -272 -1985 -255
rect -1885 -255 -1835 -238
rect -1777 -238 -1577 -200
rect -1777 -255 -1727 -238
rect -1885 -272 -1869 -255
rect -2001 -288 -1869 -272
rect -1743 -272 -1727 -255
rect -1627 -255 -1577 -238
rect -1519 -238 -1319 -200
rect -1519 -255 -1469 -238
rect -1627 -272 -1611 -255
rect -1743 -288 -1611 -272
rect -1485 -272 -1469 -255
rect -1369 -255 -1319 -238
rect -1261 -238 -1061 -200
rect -1261 -255 -1211 -238
rect -1369 -272 -1353 -255
rect -1485 -288 -1353 -272
rect -1227 -272 -1211 -255
rect -1111 -255 -1061 -238
rect -1003 -238 -803 -200
rect -1003 -255 -953 -238
rect -1111 -272 -1095 -255
rect -1227 -288 -1095 -272
rect -969 -272 -953 -255
rect -853 -255 -803 -238
rect -745 -238 -545 -200
rect -745 -255 -695 -238
rect -853 -272 -837 -255
rect -969 -288 -837 -272
rect -711 -272 -695 -255
rect -595 -255 -545 -238
rect -487 -238 -287 -200
rect -487 -255 -437 -238
rect -595 -272 -579 -255
rect -711 -288 -579 -272
rect -453 -272 -437 -255
rect -337 -255 -287 -238
rect -229 -238 -29 -200
rect -229 -255 -179 -238
rect -337 -272 -321 -255
rect -453 -288 -321 -272
rect -195 -272 -179 -255
rect -79 -255 -29 -238
rect 29 -238 229 -200
rect 29 -255 79 -238
rect -79 -272 -63 -255
rect -195 -288 -63 -272
rect 63 -272 79 -255
rect 179 -255 229 -238
rect 287 -238 487 -200
rect 287 -255 337 -238
rect 179 -272 195 -255
rect 63 -288 195 -272
rect 321 -272 337 -255
rect 437 -255 487 -238
rect 545 -238 745 -200
rect 545 -255 595 -238
rect 437 -272 453 -255
rect 321 -288 453 -272
rect 579 -272 595 -255
rect 695 -255 745 -238
rect 803 -238 1003 -200
rect 803 -255 853 -238
rect 695 -272 711 -255
rect 579 -288 711 -272
rect 837 -272 853 -255
rect 953 -255 1003 -238
rect 1061 -238 1261 -200
rect 1061 -255 1111 -238
rect 953 -272 969 -255
rect 837 -288 969 -272
rect 1095 -272 1111 -255
rect 1211 -255 1261 -238
rect 1319 -238 1519 -200
rect 1319 -255 1369 -238
rect 1211 -272 1227 -255
rect 1095 -288 1227 -272
rect 1353 -272 1369 -255
rect 1469 -255 1519 -238
rect 1577 -238 1777 -200
rect 1577 -255 1627 -238
rect 1469 -272 1485 -255
rect 1353 -288 1485 -272
rect 1611 -272 1627 -255
rect 1727 -255 1777 -238
rect 1835 -238 2035 -200
rect 1835 -255 1885 -238
rect 1727 -272 1743 -255
rect 1611 -288 1743 -272
rect 1869 -272 1885 -255
rect 1985 -255 2035 -238
rect 2093 -238 2293 -200
rect 2093 -255 2143 -238
rect 1985 -272 2001 -255
rect 1869 -288 2001 -272
rect 2127 -272 2143 -255
rect 2243 -255 2293 -238
rect 2351 -238 2551 -200
rect 2351 -255 2401 -238
rect 2243 -272 2259 -255
rect 2127 -288 2259 -272
rect 2385 -272 2401 -255
rect 2501 -255 2551 -238
rect 2609 -238 2809 -200
rect 2609 -255 2659 -238
rect 2501 -272 2517 -255
rect 2385 -288 2517 -272
rect 2643 -272 2659 -255
rect 2759 -255 2809 -238
rect 2867 -238 3067 -200
rect 2867 -255 2917 -238
rect 2759 -272 2775 -255
rect 2643 -288 2775 -272
rect 2901 -272 2917 -255
rect 3017 -255 3067 -238
rect 3125 -238 3325 -200
rect 3125 -255 3175 -238
rect 3017 -272 3033 -255
rect 2901 -288 3033 -272
rect 3159 -272 3175 -255
rect 3275 -255 3325 -238
rect 3383 -238 3583 -200
rect 3383 -255 3433 -238
rect 3275 -272 3291 -255
rect 3159 -288 3291 -272
rect 3417 -272 3433 -255
rect 3533 -255 3583 -238
rect 3641 -238 3841 -200
rect 3641 -255 3691 -238
rect 3533 -272 3549 -255
rect 3417 -288 3549 -272
rect 3675 -272 3691 -255
rect 3791 -255 3841 -238
rect 3899 -238 4099 -200
rect 3899 -255 3949 -238
rect 3791 -272 3807 -255
rect 3675 -288 3807 -272
rect 3933 -272 3949 -255
rect 4049 -255 4099 -238
rect 4157 -238 4357 -200
rect 4157 -255 4207 -238
rect 4049 -272 4065 -255
rect 3933 -288 4065 -272
rect 4191 -272 4207 -255
rect 4307 -255 4357 -238
rect 4415 -238 4615 -200
rect 4415 -255 4465 -238
rect 4307 -272 4323 -255
rect 4191 -288 4323 -272
rect 4449 -272 4465 -255
rect 4565 -255 4615 -238
rect 4673 -238 4873 -200
rect 4673 -255 4723 -238
rect 4565 -272 4581 -255
rect 4449 -288 4581 -272
rect 4707 -272 4723 -255
rect 4823 -255 4873 -238
rect 4931 -238 5131 -200
rect 4931 -255 4981 -238
rect 4823 -272 4839 -255
rect 4707 -288 4839 -272
rect 4965 -272 4981 -255
rect 5081 -255 5131 -238
rect 5081 -272 5097 -255
rect 4965 -288 5097 -272
<< polycont >>
rect -5081 238 -4981 272
rect -4823 238 -4723 272
rect -4565 238 -4465 272
rect -4307 238 -4207 272
rect -4049 238 -3949 272
rect -3791 238 -3691 272
rect -3533 238 -3433 272
rect -3275 238 -3175 272
rect -3017 238 -2917 272
rect -2759 238 -2659 272
rect -2501 238 -2401 272
rect -2243 238 -2143 272
rect -1985 238 -1885 272
rect -1727 238 -1627 272
rect -1469 238 -1369 272
rect -1211 238 -1111 272
rect -953 238 -853 272
rect -695 238 -595 272
rect -437 238 -337 272
rect -179 238 -79 272
rect 79 238 179 272
rect 337 238 437 272
rect 595 238 695 272
rect 853 238 953 272
rect 1111 238 1211 272
rect 1369 238 1469 272
rect 1627 238 1727 272
rect 1885 238 1985 272
rect 2143 238 2243 272
rect 2401 238 2501 272
rect 2659 238 2759 272
rect 2917 238 3017 272
rect 3175 238 3275 272
rect 3433 238 3533 272
rect 3691 238 3791 272
rect 3949 238 4049 272
rect 4207 238 4307 272
rect 4465 238 4565 272
rect 4723 238 4823 272
rect 4981 238 5081 272
rect -5081 -272 -4981 -238
rect -4823 -272 -4723 -238
rect -4565 -272 -4465 -238
rect -4307 -272 -4207 -238
rect -4049 -272 -3949 -238
rect -3791 -272 -3691 -238
rect -3533 -272 -3433 -238
rect -3275 -272 -3175 -238
rect -3017 -272 -2917 -238
rect -2759 -272 -2659 -238
rect -2501 -272 -2401 -238
rect -2243 -272 -2143 -238
rect -1985 -272 -1885 -238
rect -1727 -272 -1627 -238
rect -1469 -272 -1369 -238
rect -1211 -272 -1111 -238
rect -953 -272 -853 -238
rect -695 -272 -595 -238
rect -437 -272 -337 -238
rect -179 -272 -79 -238
rect 79 -272 179 -238
rect 337 -272 437 -238
rect 595 -272 695 -238
rect 853 -272 953 -238
rect 1111 -272 1211 -238
rect 1369 -272 1469 -238
rect 1627 -272 1727 -238
rect 1885 -272 1985 -238
rect 2143 -272 2243 -238
rect 2401 -272 2501 -238
rect 2659 -272 2759 -238
rect 2917 -272 3017 -238
rect 3175 -272 3275 -238
rect 3433 -272 3533 -238
rect 3691 -272 3791 -238
rect 3949 -272 4049 -238
rect 4207 -272 4307 -238
rect 4465 -272 4565 -238
rect 4723 -272 4823 -238
rect 4981 -272 5081 -238
<< locali >>
rect -5311 376 -5215 410
rect 5215 376 5311 410
rect -5311 314 -5277 376
rect 5277 314 5311 376
rect -5097 238 -5081 272
rect -4981 238 -4965 272
rect -4839 238 -4823 272
rect -4723 238 -4707 272
rect -4581 238 -4565 272
rect -4465 238 -4449 272
rect -4323 238 -4307 272
rect -4207 238 -4191 272
rect -4065 238 -4049 272
rect -3949 238 -3933 272
rect -3807 238 -3791 272
rect -3691 238 -3675 272
rect -3549 238 -3533 272
rect -3433 238 -3417 272
rect -3291 238 -3275 272
rect -3175 238 -3159 272
rect -3033 238 -3017 272
rect -2917 238 -2901 272
rect -2775 238 -2759 272
rect -2659 238 -2643 272
rect -2517 238 -2501 272
rect -2401 238 -2385 272
rect -2259 238 -2243 272
rect -2143 238 -2127 272
rect -2001 238 -1985 272
rect -1885 238 -1869 272
rect -1743 238 -1727 272
rect -1627 238 -1611 272
rect -1485 238 -1469 272
rect -1369 238 -1353 272
rect -1227 238 -1211 272
rect -1111 238 -1095 272
rect -969 238 -953 272
rect -853 238 -837 272
rect -711 238 -695 272
rect -595 238 -579 272
rect -453 238 -437 272
rect -337 238 -321 272
rect -195 238 -179 272
rect -79 238 -63 272
rect 63 238 79 272
rect 179 238 195 272
rect 321 238 337 272
rect 437 238 453 272
rect 579 238 595 272
rect 695 238 711 272
rect 837 238 853 272
rect 953 238 969 272
rect 1095 238 1111 272
rect 1211 238 1227 272
rect 1353 238 1369 272
rect 1469 238 1485 272
rect 1611 238 1627 272
rect 1727 238 1743 272
rect 1869 238 1885 272
rect 1985 238 2001 272
rect 2127 238 2143 272
rect 2243 238 2259 272
rect 2385 238 2401 272
rect 2501 238 2517 272
rect 2643 238 2659 272
rect 2759 238 2775 272
rect 2901 238 2917 272
rect 3017 238 3033 272
rect 3159 238 3175 272
rect 3275 238 3291 272
rect 3417 238 3433 272
rect 3533 238 3549 272
rect 3675 238 3691 272
rect 3791 238 3807 272
rect 3933 238 3949 272
rect 4049 238 4065 272
rect 4191 238 4207 272
rect 4307 238 4323 272
rect 4449 238 4465 272
rect 4565 238 4581 272
rect 4707 238 4723 272
rect 4823 238 4839 272
rect 4965 238 4981 272
rect 5081 238 5097 272
rect -5177 188 -5143 204
rect -5177 -204 -5143 -188
rect -4919 188 -4885 204
rect -4919 -204 -4885 -188
rect -4661 188 -4627 204
rect -4661 -204 -4627 -188
rect -4403 188 -4369 204
rect -4403 -204 -4369 -188
rect -4145 188 -4111 204
rect -4145 -204 -4111 -188
rect -3887 188 -3853 204
rect -3887 -204 -3853 -188
rect -3629 188 -3595 204
rect -3629 -204 -3595 -188
rect -3371 188 -3337 204
rect -3371 -204 -3337 -188
rect -3113 188 -3079 204
rect -3113 -204 -3079 -188
rect -2855 188 -2821 204
rect -2855 -204 -2821 -188
rect -2597 188 -2563 204
rect -2597 -204 -2563 -188
rect -2339 188 -2305 204
rect -2339 -204 -2305 -188
rect -2081 188 -2047 204
rect -2081 -204 -2047 -188
rect -1823 188 -1789 204
rect -1823 -204 -1789 -188
rect -1565 188 -1531 204
rect -1565 -204 -1531 -188
rect -1307 188 -1273 204
rect -1307 -204 -1273 -188
rect -1049 188 -1015 204
rect -1049 -204 -1015 -188
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect 1015 188 1049 204
rect 1015 -204 1049 -188
rect 1273 188 1307 204
rect 1273 -204 1307 -188
rect 1531 188 1565 204
rect 1531 -204 1565 -188
rect 1789 188 1823 204
rect 1789 -204 1823 -188
rect 2047 188 2081 204
rect 2047 -204 2081 -188
rect 2305 188 2339 204
rect 2305 -204 2339 -188
rect 2563 188 2597 204
rect 2563 -204 2597 -188
rect 2821 188 2855 204
rect 2821 -204 2855 -188
rect 3079 188 3113 204
rect 3079 -204 3113 -188
rect 3337 188 3371 204
rect 3337 -204 3371 -188
rect 3595 188 3629 204
rect 3595 -204 3629 -188
rect 3853 188 3887 204
rect 3853 -204 3887 -188
rect 4111 188 4145 204
rect 4111 -204 4145 -188
rect 4369 188 4403 204
rect 4369 -204 4403 -188
rect 4627 188 4661 204
rect 4627 -204 4661 -188
rect 4885 188 4919 204
rect 4885 -204 4919 -188
rect 5143 188 5177 204
rect 5143 -204 5177 -188
rect -5097 -272 -5081 -238
rect -4981 -272 -4965 -238
rect -4839 -272 -4823 -238
rect -4723 -272 -4707 -238
rect -4581 -272 -4565 -238
rect -4465 -272 -4449 -238
rect -4323 -272 -4307 -238
rect -4207 -272 -4191 -238
rect -4065 -272 -4049 -238
rect -3949 -272 -3933 -238
rect -3807 -272 -3791 -238
rect -3691 -272 -3675 -238
rect -3549 -272 -3533 -238
rect -3433 -272 -3417 -238
rect -3291 -272 -3275 -238
rect -3175 -272 -3159 -238
rect -3033 -272 -3017 -238
rect -2917 -272 -2901 -238
rect -2775 -272 -2759 -238
rect -2659 -272 -2643 -238
rect -2517 -272 -2501 -238
rect -2401 -272 -2385 -238
rect -2259 -272 -2243 -238
rect -2143 -272 -2127 -238
rect -2001 -272 -1985 -238
rect -1885 -272 -1869 -238
rect -1743 -272 -1727 -238
rect -1627 -272 -1611 -238
rect -1485 -272 -1469 -238
rect -1369 -272 -1353 -238
rect -1227 -272 -1211 -238
rect -1111 -272 -1095 -238
rect -969 -272 -953 -238
rect -853 -272 -837 -238
rect -711 -272 -695 -238
rect -595 -272 -579 -238
rect -453 -272 -437 -238
rect -337 -272 -321 -238
rect -195 -272 -179 -238
rect -79 -272 -63 -238
rect 63 -272 79 -238
rect 179 -272 195 -238
rect 321 -272 337 -238
rect 437 -272 453 -238
rect 579 -272 595 -238
rect 695 -272 711 -238
rect 837 -272 853 -238
rect 953 -272 969 -238
rect 1095 -272 1111 -238
rect 1211 -272 1227 -238
rect 1353 -272 1369 -238
rect 1469 -272 1485 -238
rect 1611 -272 1627 -238
rect 1727 -272 1743 -238
rect 1869 -272 1885 -238
rect 1985 -272 2001 -238
rect 2127 -272 2143 -238
rect 2243 -272 2259 -238
rect 2385 -272 2401 -238
rect 2501 -272 2517 -238
rect 2643 -272 2659 -238
rect 2759 -272 2775 -238
rect 2901 -272 2917 -238
rect 3017 -272 3033 -238
rect 3159 -272 3175 -238
rect 3275 -272 3291 -238
rect 3417 -272 3433 -238
rect 3533 -272 3549 -238
rect 3675 -272 3691 -238
rect 3791 -272 3807 -238
rect 3933 -272 3949 -238
rect 4049 -272 4065 -238
rect 4191 -272 4207 -238
rect 4307 -272 4323 -238
rect 4449 -272 4465 -238
rect 4565 -272 4581 -238
rect 4707 -272 4723 -238
rect 4823 -272 4839 -238
rect 4965 -272 4981 -238
rect 5081 -272 5097 -238
rect -5311 -376 -5277 -314
rect 5277 -376 5311 -314
rect -5311 -410 -5215 -376
rect 5215 -410 5311 -376
<< viali >>
rect -5081 238 -4981 272
rect -4823 238 -4723 272
rect -4565 238 -4465 272
rect -4307 238 -4207 272
rect -4049 238 -3949 272
rect -3791 238 -3691 272
rect -3533 238 -3433 272
rect -3275 238 -3175 272
rect -3017 238 -2917 272
rect -2759 238 -2659 272
rect -2501 238 -2401 272
rect -2243 238 -2143 272
rect -1985 238 -1885 272
rect -1727 238 -1627 272
rect -1469 238 -1369 272
rect -1211 238 -1111 272
rect -953 238 -853 272
rect -695 238 -595 272
rect -437 238 -337 272
rect -179 238 -79 272
rect 79 238 179 272
rect 337 238 437 272
rect 595 238 695 272
rect 853 238 953 272
rect 1111 238 1211 272
rect 1369 238 1469 272
rect 1627 238 1727 272
rect 1885 238 1985 272
rect 2143 238 2243 272
rect 2401 238 2501 272
rect 2659 238 2759 272
rect 2917 238 3017 272
rect 3175 238 3275 272
rect 3433 238 3533 272
rect 3691 238 3791 272
rect 3949 238 4049 272
rect 4207 238 4307 272
rect 4465 238 4565 272
rect 4723 238 4823 272
rect 4981 238 5081 272
rect -5177 -188 -5143 188
rect -4919 -188 -4885 188
rect -4661 -188 -4627 188
rect -4403 -188 -4369 188
rect -4145 -188 -4111 188
rect -3887 -188 -3853 188
rect -3629 -188 -3595 188
rect -3371 -188 -3337 188
rect -3113 -188 -3079 188
rect -2855 -188 -2821 188
rect -2597 -188 -2563 188
rect -2339 -188 -2305 188
rect -2081 -188 -2047 188
rect -1823 -188 -1789 188
rect -1565 -188 -1531 188
rect -1307 -188 -1273 188
rect -1049 -188 -1015 188
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect 1015 -188 1049 188
rect 1273 -188 1307 188
rect 1531 -188 1565 188
rect 1789 -188 1823 188
rect 2047 -188 2081 188
rect 2305 -188 2339 188
rect 2563 -188 2597 188
rect 2821 -188 2855 188
rect 3079 -188 3113 188
rect 3337 -188 3371 188
rect 3595 -188 3629 188
rect 3853 -188 3887 188
rect 4111 -188 4145 188
rect 4369 -188 4403 188
rect 4627 -188 4661 188
rect 4885 -188 4919 188
rect 5143 -188 5177 188
rect -5081 -272 -4981 -238
rect -4823 -272 -4723 -238
rect -4565 -272 -4465 -238
rect -4307 -272 -4207 -238
rect -4049 -272 -3949 -238
rect -3791 -272 -3691 -238
rect -3533 -272 -3433 -238
rect -3275 -272 -3175 -238
rect -3017 -272 -2917 -238
rect -2759 -272 -2659 -238
rect -2501 -272 -2401 -238
rect -2243 -272 -2143 -238
rect -1985 -272 -1885 -238
rect -1727 -272 -1627 -238
rect -1469 -272 -1369 -238
rect -1211 -272 -1111 -238
rect -953 -272 -853 -238
rect -695 -272 -595 -238
rect -437 -272 -337 -238
rect -179 -272 -79 -238
rect 79 -272 179 -238
rect 337 -272 437 -238
rect 595 -272 695 -238
rect 853 -272 953 -238
rect 1111 -272 1211 -238
rect 1369 -272 1469 -238
rect 1627 -272 1727 -238
rect 1885 -272 1985 -238
rect 2143 -272 2243 -238
rect 2401 -272 2501 -238
rect 2659 -272 2759 -238
rect 2917 -272 3017 -238
rect 3175 -272 3275 -238
rect 3433 -272 3533 -238
rect 3691 -272 3791 -238
rect 3949 -272 4049 -238
rect 4207 -272 4307 -238
rect 4465 -272 4565 -238
rect 4723 -272 4823 -238
rect 4981 -272 5081 -238
<< metal1 >>
rect -5093 272 -4969 278
rect -5093 238 -5081 272
rect -4981 238 -4969 272
rect -5093 232 -4969 238
rect -4835 272 -4711 278
rect -4835 238 -4823 272
rect -4723 238 -4711 272
rect -4835 232 -4711 238
rect -4577 272 -4453 278
rect -4577 238 -4565 272
rect -4465 238 -4453 272
rect -4577 232 -4453 238
rect -4319 272 -4195 278
rect -4319 238 -4307 272
rect -4207 238 -4195 272
rect -4319 232 -4195 238
rect -4061 272 -3937 278
rect -4061 238 -4049 272
rect -3949 238 -3937 272
rect -4061 232 -3937 238
rect -3803 272 -3679 278
rect -3803 238 -3791 272
rect -3691 238 -3679 272
rect -3803 232 -3679 238
rect -3545 272 -3421 278
rect -3545 238 -3533 272
rect -3433 238 -3421 272
rect -3545 232 -3421 238
rect -3287 272 -3163 278
rect -3287 238 -3275 272
rect -3175 238 -3163 272
rect -3287 232 -3163 238
rect -3029 272 -2905 278
rect -3029 238 -3017 272
rect -2917 238 -2905 272
rect -3029 232 -2905 238
rect -2771 272 -2647 278
rect -2771 238 -2759 272
rect -2659 238 -2647 272
rect -2771 232 -2647 238
rect -2513 272 -2389 278
rect -2513 238 -2501 272
rect -2401 238 -2389 272
rect -2513 232 -2389 238
rect -2255 272 -2131 278
rect -2255 238 -2243 272
rect -2143 238 -2131 272
rect -2255 232 -2131 238
rect -1997 272 -1873 278
rect -1997 238 -1985 272
rect -1885 238 -1873 272
rect -1997 232 -1873 238
rect -1739 272 -1615 278
rect -1739 238 -1727 272
rect -1627 238 -1615 272
rect -1739 232 -1615 238
rect -1481 272 -1357 278
rect -1481 238 -1469 272
rect -1369 238 -1357 272
rect -1481 232 -1357 238
rect -1223 272 -1099 278
rect -1223 238 -1211 272
rect -1111 238 -1099 272
rect -1223 232 -1099 238
rect -965 272 -841 278
rect -965 238 -953 272
rect -853 238 -841 272
rect -965 232 -841 238
rect -707 272 -583 278
rect -707 238 -695 272
rect -595 238 -583 272
rect -707 232 -583 238
rect -449 272 -325 278
rect -449 238 -437 272
rect -337 238 -325 272
rect -449 232 -325 238
rect -191 272 -67 278
rect -191 238 -179 272
rect -79 238 -67 272
rect -191 232 -67 238
rect 67 272 191 278
rect 67 238 79 272
rect 179 238 191 272
rect 67 232 191 238
rect 325 272 449 278
rect 325 238 337 272
rect 437 238 449 272
rect 325 232 449 238
rect 583 272 707 278
rect 583 238 595 272
rect 695 238 707 272
rect 583 232 707 238
rect 841 272 965 278
rect 841 238 853 272
rect 953 238 965 272
rect 841 232 965 238
rect 1099 272 1223 278
rect 1099 238 1111 272
rect 1211 238 1223 272
rect 1099 232 1223 238
rect 1357 272 1481 278
rect 1357 238 1369 272
rect 1469 238 1481 272
rect 1357 232 1481 238
rect 1615 272 1739 278
rect 1615 238 1627 272
rect 1727 238 1739 272
rect 1615 232 1739 238
rect 1873 272 1997 278
rect 1873 238 1885 272
rect 1985 238 1997 272
rect 1873 232 1997 238
rect 2131 272 2255 278
rect 2131 238 2143 272
rect 2243 238 2255 272
rect 2131 232 2255 238
rect 2389 272 2513 278
rect 2389 238 2401 272
rect 2501 238 2513 272
rect 2389 232 2513 238
rect 2647 272 2771 278
rect 2647 238 2659 272
rect 2759 238 2771 272
rect 2647 232 2771 238
rect 2905 272 3029 278
rect 2905 238 2917 272
rect 3017 238 3029 272
rect 2905 232 3029 238
rect 3163 272 3287 278
rect 3163 238 3175 272
rect 3275 238 3287 272
rect 3163 232 3287 238
rect 3421 272 3545 278
rect 3421 238 3433 272
rect 3533 238 3545 272
rect 3421 232 3545 238
rect 3679 272 3803 278
rect 3679 238 3691 272
rect 3791 238 3803 272
rect 3679 232 3803 238
rect 3937 272 4061 278
rect 3937 238 3949 272
rect 4049 238 4061 272
rect 3937 232 4061 238
rect 4195 272 4319 278
rect 4195 238 4207 272
rect 4307 238 4319 272
rect 4195 232 4319 238
rect 4453 272 4577 278
rect 4453 238 4465 272
rect 4565 238 4577 272
rect 4453 232 4577 238
rect 4711 272 4835 278
rect 4711 238 4723 272
rect 4823 238 4835 272
rect 4711 232 4835 238
rect 4969 272 5093 278
rect 4969 238 4981 272
rect 5081 238 5093 272
rect 4969 232 5093 238
rect -5183 188 -5137 200
rect -5183 -188 -5177 188
rect -5143 -188 -5137 188
rect -5183 -200 -5137 -188
rect -4925 188 -4879 200
rect -4925 -188 -4919 188
rect -4885 -188 -4879 188
rect -4925 -200 -4879 -188
rect -4667 188 -4621 200
rect -4667 -188 -4661 188
rect -4627 -188 -4621 188
rect -4667 -200 -4621 -188
rect -4409 188 -4363 200
rect -4409 -188 -4403 188
rect -4369 -188 -4363 188
rect -4409 -200 -4363 -188
rect -4151 188 -4105 200
rect -4151 -188 -4145 188
rect -4111 -188 -4105 188
rect -4151 -200 -4105 -188
rect -3893 188 -3847 200
rect -3893 -188 -3887 188
rect -3853 -188 -3847 188
rect -3893 -200 -3847 -188
rect -3635 188 -3589 200
rect -3635 -188 -3629 188
rect -3595 -188 -3589 188
rect -3635 -200 -3589 -188
rect -3377 188 -3331 200
rect -3377 -188 -3371 188
rect -3337 -188 -3331 188
rect -3377 -200 -3331 -188
rect -3119 188 -3073 200
rect -3119 -188 -3113 188
rect -3079 -188 -3073 188
rect -3119 -200 -3073 -188
rect -2861 188 -2815 200
rect -2861 -188 -2855 188
rect -2821 -188 -2815 188
rect -2861 -200 -2815 -188
rect -2603 188 -2557 200
rect -2603 -188 -2597 188
rect -2563 -188 -2557 188
rect -2603 -200 -2557 -188
rect -2345 188 -2299 200
rect -2345 -188 -2339 188
rect -2305 -188 -2299 188
rect -2345 -200 -2299 -188
rect -2087 188 -2041 200
rect -2087 -188 -2081 188
rect -2047 -188 -2041 188
rect -2087 -200 -2041 -188
rect -1829 188 -1783 200
rect -1829 -188 -1823 188
rect -1789 -188 -1783 188
rect -1829 -200 -1783 -188
rect -1571 188 -1525 200
rect -1571 -188 -1565 188
rect -1531 -188 -1525 188
rect -1571 -200 -1525 -188
rect -1313 188 -1267 200
rect -1313 -188 -1307 188
rect -1273 -188 -1267 188
rect -1313 -200 -1267 -188
rect -1055 188 -1009 200
rect -1055 -188 -1049 188
rect -1015 -188 -1009 188
rect -1055 -200 -1009 -188
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect 1009 188 1055 200
rect 1009 -188 1015 188
rect 1049 -188 1055 188
rect 1009 -200 1055 -188
rect 1267 188 1313 200
rect 1267 -188 1273 188
rect 1307 -188 1313 188
rect 1267 -200 1313 -188
rect 1525 188 1571 200
rect 1525 -188 1531 188
rect 1565 -188 1571 188
rect 1525 -200 1571 -188
rect 1783 188 1829 200
rect 1783 -188 1789 188
rect 1823 -188 1829 188
rect 1783 -200 1829 -188
rect 2041 188 2087 200
rect 2041 -188 2047 188
rect 2081 -188 2087 188
rect 2041 -200 2087 -188
rect 2299 188 2345 200
rect 2299 -188 2305 188
rect 2339 -188 2345 188
rect 2299 -200 2345 -188
rect 2557 188 2603 200
rect 2557 -188 2563 188
rect 2597 -188 2603 188
rect 2557 -200 2603 -188
rect 2815 188 2861 200
rect 2815 -188 2821 188
rect 2855 -188 2861 188
rect 2815 -200 2861 -188
rect 3073 188 3119 200
rect 3073 -188 3079 188
rect 3113 -188 3119 188
rect 3073 -200 3119 -188
rect 3331 188 3377 200
rect 3331 -188 3337 188
rect 3371 -188 3377 188
rect 3331 -200 3377 -188
rect 3589 188 3635 200
rect 3589 -188 3595 188
rect 3629 -188 3635 188
rect 3589 -200 3635 -188
rect 3847 188 3893 200
rect 3847 -188 3853 188
rect 3887 -188 3893 188
rect 3847 -200 3893 -188
rect 4105 188 4151 200
rect 4105 -188 4111 188
rect 4145 -188 4151 188
rect 4105 -200 4151 -188
rect 4363 188 4409 200
rect 4363 -188 4369 188
rect 4403 -188 4409 188
rect 4363 -200 4409 -188
rect 4621 188 4667 200
rect 4621 -188 4627 188
rect 4661 -188 4667 188
rect 4621 -200 4667 -188
rect 4879 188 4925 200
rect 4879 -188 4885 188
rect 4919 -188 4925 188
rect 4879 -200 4925 -188
rect 5137 188 5183 200
rect 5137 -188 5143 188
rect 5177 -188 5183 188
rect 5137 -200 5183 -188
rect -5093 -238 -4969 -232
rect -5093 -272 -5081 -238
rect -4981 -272 -4969 -238
rect -5093 -278 -4969 -272
rect -4835 -238 -4711 -232
rect -4835 -272 -4823 -238
rect -4723 -272 -4711 -238
rect -4835 -278 -4711 -272
rect -4577 -238 -4453 -232
rect -4577 -272 -4565 -238
rect -4465 -272 -4453 -238
rect -4577 -278 -4453 -272
rect -4319 -238 -4195 -232
rect -4319 -272 -4307 -238
rect -4207 -272 -4195 -238
rect -4319 -278 -4195 -272
rect -4061 -238 -3937 -232
rect -4061 -272 -4049 -238
rect -3949 -272 -3937 -238
rect -4061 -278 -3937 -272
rect -3803 -238 -3679 -232
rect -3803 -272 -3791 -238
rect -3691 -272 -3679 -238
rect -3803 -278 -3679 -272
rect -3545 -238 -3421 -232
rect -3545 -272 -3533 -238
rect -3433 -272 -3421 -238
rect -3545 -278 -3421 -272
rect -3287 -238 -3163 -232
rect -3287 -272 -3275 -238
rect -3175 -272 -3163 -238
rect -3287 -278 -3163 -272
rect -3029 -238 -2905 -232
rect -3029 -272 -3017 -238
rect -2917 -272 -2905 -238
rect -3029 -278 -2905 -272
rect -2771 -238 -2647 -232
rect -2771 -272 -2759 -238
rect -2659 -272 -2647 -238
rect -2771 -278 -2647 -272
rect -2513 -238 -2389 -232
rect -2513 -272 -2501 -238
rect -2401 -272 -2389 -238
rect -2513 -278 -2389 -272
rect -2255 -238 -2131 -232
rect -2255 -272 -2243 -238
rect -2143 -272 -2131 -238
rect -2255 -278 -2131 -272
rect -1997 -238 -1873 -232
rect -1997 -272 -1985 -238
rect -1885 -272 -1873 -238
rect -1997 -278 -1873 -272
rect -1739 -238 -1615 -232
rect -1739 -272 -1727 -238
rect -1627 -272 -1615 -238
rect -1739 -278 -1615 -272
rect -1481 -238 -1357 -232
rect -1481 -272 -1469 -238
rect -1369 -272 -1357 -238
rect -1481 -278 -1357 -272
rect -1223 -238 -1099 -232
rect -1223 -272 -1211 -238
rect -1111 -272 -1099 -238
rect -1223 -278 -1099 -272
rect -965 -238 -841 -232
rect -965 -272 -953 -238
rect -853 -272 -841 -238
rect -965 -278 -841 -272
rect -707 -238 -583 -232
rect -707 -272 -695 -238
rect -595 -272 -583 -238
rect -707 -278 -583 -272
rect -449 -238 -325 -232
rect -449 -272 -437 -238
rect -337 -272 -325 -238
rect -449 -278 -325 -272
rect -191 -238 -67 -232
rect -191 -272 -179 -238
rect -79 -272 -67 -238
rect -191 -278 -67 -272
rect 67 -238 191 -232
rect 67 -272 79 -238
rect 179 -272 191 -238
rect 67 -278 191 -272
rect 325 -238 449 -232
rect 325 -272 337 -238
rect 437 -272 449 -238
rect 325 -278 449 -272
rect 583 -238 707 -232
rect 583 -272 595 -238
rect 695 -272 707 -238
rect 583 -278 707 -272
rect 841 -238 965 -232
rect 841 -272 853 -238
rect 953 -272 965 -238
rect 841 -278 965 -272
rect 1099 -238 1223 -232
rect 1099 -272 1111 -238
rect 1211 -272 1223 -238
rect 1099 -278 1223 -272
rect 1357 -238 1481 -232
rect 1357 -272 1369 -238
rect 1469 -272 1481 -238
rect 1357 -278 1481 -272
rect 1615 -238 1739 -232
rect 1615 -272 1627 -238
rect 1727 -272 1739 -238
rect 1615 -278 1739 -272
rect 1873 -238 1997 -232
rect 1873 -272 1885 -238
rect 1985 -272 1997 -238
rect 1873 -278 1997 -272
rect 2131 -238 2255 -232
rect 2131 -272 2143 -238
rect 2243 -272 2255 -238
rect 2131 -278 2255 -272
rect 2389 -238 2513 -232
rect 2389 -272 2401 -238
rect 2501 -272 2513 -238
rect 2389 -278 2513 -272
rect 2647 -238 2771 -232
rect 2647 -272 2659 -238
rect 2759 -272 2771 -238
rect 2647 -278 2771 -272
rect 2905 -238 3029 -232
rect 2905 -272 2917 -238
rect 3017 -272 3029 -238
rect 2905 -278 3029 -272
rect 3163 -238 3287 -232
rect 3163 -272 3175 -238
rect 3275 -272 3287 -238
rect 3163 -278 3287 -272
rect 3421 -238 3545 -232
rect 3421 -272 3433 -238
rect 3533 -272 3545 -238
rect 3421 -278 3545 -272
rect 3679 -238 3803 -232
rect 3679 -272 3691 -238
rect 3791 -272 3803 -238
rect 3679 -278 3803 -272
rect 3937 -238 4061 -232
rect 3937 -272 3949 -238
rect 4049 -272 4061 -238
rect 3937 -278 4061 -272
rect 4195 -238 4319 -232
rect 4195 -272 4207 -238
rect 4307 -272 4319 -238
rect 4195 -278 4319 -272
rect 4453 -238 4577 -232
rect 4453 -272 4465 -238
rect 4565 -272 4577 -238
rect 4453 -278 4577 -272
rect 4711 -238 4835 -232
rect 4711 -272 4723 -238
rect 4823 -272 4835 -238
rect 4711 -278 4835 -272
rect 4969 -238 5093 -232
rect 4969 -272 4981 -238
rect 5081 -272 5093 -238
rect 4969 -278 5093 -272
<< properties >>
string FIXED_BBOX -5294 -393 5294 393
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2 l 1 m 1 nf 40 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

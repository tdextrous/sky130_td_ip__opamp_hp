magic
tech sky130A
magscale 1 2
timestamp 1713394428
<< nwell >>
rect -3067 -1197 3067 1197
<< mvpmos >>
rect -2809 -900 -2609 900
rect -2551 -900 -2351 900
rect -2293 -900 -2093 900
rect -2035 -900 -1835 900
rect -1777 -900 -1577 900
rect -1519 -900 -1319 900
rect -1261 -900 -1061 900
rect -1003 -900 -803 900
rect -745 -900 -545 900
rect -487 -900 -287 900
rect -229 -900 -29 900
rect 29 -900 229 900
rect 287 -900 487 900
rect 545 -900 745 900
rect 803 -900 1003 900
rect 1061 -900 1261 900
rect 1319 -900 1519 900
rect 1577 -900 1777 900
rect 1835 -900 2035 900
rect 2093 -900 2293 900
rect 2351 -900 2551 900
rect 2609 -900 2809 900
<< mvpdiff >>
rect -2867 888 -2809 900
rect -2867 -888 -2855 888
rect -2821 -888 -2809 888
rect -2867 -900 -2809 -888
rect -2609 888 -2551 900
rect -2609 -888 -2597 888
rect -2563 -888 -2551 888
rect -2609 -900 -2551 -888
rect -2351 888 -2293 900
rect -2351 -888 -2339 888
rect -2305 -888 -2293 888
rect -2351 -900 -2293 -888
rect -2093 888 -2035 900
rect -2093 -888 -2081 888
rect -2047 -888 -2035 888
rect -2093 -900 -2035 -888
rect -1835 888 -1777 900
rect -1835 -888 -1823 888
rect -1789 -888 -1777 888
rect -1835 -900 -1777 -888
rect -1577 888 -1519 900
rect -1577 -888 -1565 888
rect -1531 -888 -1519 888
rect -1577 -900 -1519 -888
rect -1319 888 -1261 900
rect -1319 -888 -1307 888
rect -1273 -888 -1261 888
rect -1319 -900 -1261 -888
rect -1061 888 -1003 900
rect -1061 -888 -1049 888
rect -1015 -888 -1003 888
rect -1061 -900 -1003 -888
rect -803 888 -745 900
rect -803 -888 -791 888
rect -757 -888 -745 888
rect -803 -900 -745 -888
rect -545 888 -487 900
rect -545 -888 -533 888
rect -499 -888 -487 888
rect -545 -900 -487 -888
rect -287 888 -229 900
rect -287 -888 -275 888
rect -241 -888 -229 888
rect -287 -900 -229 -888
rect -29 888 29 900
rect -29 -888 -17 888
rect 17 -888 29 888
rect -29 -900 29 -888
rect 229 888 287 900
rect 229 -888 241 888
rect 275 -888 287 888
rect 229 -900 287 -888
rect 487 888 545 900
rect 487 -888 499 888
rect 533 -888 545 888
rect 487 -900 545 -888
rect 745 888 803 900
rect 745 -888 757 888
rect 791 -888 803 888
rect 745 -900 803 -888
rect 1003 888 1061 900
rect 1003 -888 1015 888
rect 1049 -888 1061 888
rect 1003 -900 1061 -888
rect 1261 888 1319 900
rect 1261 -888 1273 888
rect 1307 -888 1319 888
rect 1261 -900 1319 -888
rect 1519 888 1577 900
rect 1519 -888 1531 888
rect 1565 -888 1577 888
rect 1519 -900 1577 -888
rect 1777 888 1835 900
rect 1777 -888 1789 888
rect 1823 -888 1835 888
rect 1777 -900 1835 -888
rect 2035 888 2093 900
rect 2035 -888 2047 888
rect 2081 -888 2093 888
rect 2035 -900 2093 -888
rect 2293 888 2351 900
rect 2293 -888 2305 888
rect 2339 -888 2351 888
rect 2293 -900 2351 -888
rect 2551 888 2609 900
rect 2551 -888 2563 888
rect 2597 -888 2609 888
rect 2551 -900 2609 -888
rect 2809 888 2867 900
rect 2809 -888 2821 888
rect 2855 -888 2867 888
rect 2809 -900 2867 -888
<< mvpdiffc >>
rect -2855 -888 -2821 888
rect -2597 -888 -2563 888
rect -2339 -888 -2305 888
rect -2081 -888 -2047 888
rect -1823 -888 -1789 888
rect -1565 -888 -1531 888
rect -1307 -888 -1273 888
rect -1049 -888 -1015 888
rect -791 -888 -757 888
rect -533 -888 -499 888
rect -275 -888 -241 888
rect -17 -888 17 888
rect 241 -888 275 888
rect 499 -888 533 888
rect 757 -888 791 888
rect 1015 -888 1049 888
rect 1273 -888 1307 888
rect 1531 -888 1565 888
rect 1789 -888 1823 888
rect 2047 -888 2081 888
rect 2305 -888 2339 888
rect 2563 -888 2597 888
rect 2821 -888 2855 888
<< mvnsubdiff >>
rect -3001 1119 3001 1131
rect -3001 1085 -2893 1119
rect 2893 1085 3001 1119
rect -3001 1073 3001 1085
rect -3001 1023 -2943 1073
rect -3001 -1023 -2989 1023
rect -2955 -1023 -2943 1023
rect 2943 1023 3001 1073
rect -3001 -1073 -2943 -1023
rect 2943 -1023 2955 1023
rect 2989 -1023 3001 1023
rect 2943 -1073 3001 -1023
rect -3001 -1085 3001 -1073
rect -3001 -1119 -2893 -1085
rect 2893 -1119 3001 -1085
rect -3001 -1131 3001 -1119
<< mvnsubdiffcont >>
rect -2893 1085 2893 1119
rect -2989 -1023 -2955 1023
rect 2955 -1023 2989 1023
rect -2893 -1119 2893 -1085
<< poly >>
rect -2775 981 -2643 997
rect -2775 964 -2759 981
rect -2809 947 -2759 964
rect -2659 964 -2643 981
rect -2517 981 -2385 997
rect -2517 964 -2501 981
rect -2659 947 -2609 964
rect -2809 900 -2609 947
rect -2551 947 -2501 964
rect -2401 964 -2385 981
rect -2259 981 -2127 997
rect -2259 964 -2243 981
rect -2401 947 -2351 964
rect -2551 900 -2351 947
rect -2293 947 -2243 964
rect -2143 964 -2127 981
rect -2001 981 -1869 997
rect -2001 964 -1985 981
rect -2143 947 -2093 964
rect -2293 900 -2093 947
rect -2035 947 -1985 964
rect -1885 964 -1869 981
rect -1743 981 -1611 997
rect -1743 964 -1727 981
rect -1885 947 -1835 964
rect -2035 900 -1835 947
rect -1777 947 -1727 964
rect -1627 964 -1611 981
rect -1485 981 -1353 997
rect -1485 964 -1469 981
rect -1627 947 -1577 964
rect -1777 900 -1577 947
rect -1519 947 -1469 964
rect -1369 964 -1353 981
rect -1227 981 -1095 997
rect -1227 964 -1211 981
rect -1369 947 -1319 964
rect -1519 900 -1319 947
rect -1261 947 -1211 964
rect -1111 964 -1095 981
rect -969 981 -837 997
rect -969 964 -953 981
rect -1111 947 -1061 964
rect -1261 900 -1061 947
rect -1003 947 -953 964
rect -853 964 -837 981
rect -711 981 -579 997
rect -711 964 -695 981
rect -853 947 -803 964
rect -1003 900 -803 947
rect -745 947 -695 964
rect -595 964 -579 981
rect -453 981 -321 997
rect -453 964 -437 981
rect -595 947 -545 964
rect -745 900 -545 947
rect -487 947 -437 964
rect -337 964 -321 981
rect -195 981 -63 997
rect -195 964 -179 981
rect -337 947 -287 964
rect -487 900 -287 947
rect -229 947 -179 964
rect -79 964 -63 981
rect 63 981 195 997
rect 63 964 79 981
rect -79 947 -29 964
rect -229 900 -29 947
rect 29 947 79 964
rect 179 964 195 981
rect 321 981 453 997
rect 321 964 337 981
rect 179 947 229 964
rect 29 900 229 947
rect 287 947 337 964
rect 437 964 453 981
rect 579 981 711 997
rect 579 964 595 981
rect 437 947 487 964
rect 287 900 487 947
rect 545 947 595 964
rect 695 964 711 981
rect 837 981 969 997
rect 837 964 853 981
rect 695 947 745 964
rect 545 900 745 947
rect 803 947 853 964
rect 953 964 969 981
rect 1095 981 1227 997
rect 1095 964 1111 981
rect 953 947 1003 964
rect 803 900 1003 947
rect 1061 947 1111 964
rect 1211 964 1227 981
rect 1353 981 1485 997
rect 1353 964 1369 981
rect 1211 947 1261 964
rect 1061 900 1261 947
rect 1319 947 1369 964
rect 1469 964 1485 981
rect 1611 981 1743 997
rect 1611 964 1627 981
rect 1469 947 1519 964
rect 1319 900 1519 947
rect 1577 947 1627 964
rect 1727 964 1743 981
rect 1869 981 2001 997
rect 1869 964 1885 981
rect 1727 947 1777 964
rect 1577 900 1777 947
rect 1835 947 1885 964
rect 1985 964 2001 981
rect 2127 981 2259 997
rect 2127 964 2143 981
rect 1985 947 2035 964
rect 1835 900 2035 947
rect 2093 947 2143 964
rect 2243 964 2259 981
rect 2385 981 2517 997
rect 2385 964 2401 981
rect 2243 947 2293 964
rect 2093 900 2293 947
rect 2351 947 2401 964
rect 2501 964 2517 981
rect 2643 981 2775 997
rect 2643 964 2659 981
rect 2501 947 2551 964
rect 2351 900 2551 947
rect 2609 947 2659 964
rect 2759 964 2775 981
rect 2759 947 2809 964
rect 2609 900 2809 947
rect -2809 -947 -2609 -900
rect -2809 -964 -2759 -947
rect -2775 -981 -2759 -964
rect -2659 -964 -2609 -947
rect -2551 -947 -2351 -900
rect -2551 -964 -2501 -947
rect -2659 -981 -2643 -964
rect -2775 -997 -2643 -981
rect -2517 -981 -2501 -964
rect -2401 -964 -2351 -947
rect -2293 -947 -2093 -900
rect -2293 -964 -2243 -947
rect -2401 -981 -2385 -964
rect -2517 -997 -2385 -981
rect -2259 -981 -2243 -964
rect -2143 -964 -2093 -947
rect -2035 -947 -1835 -900
rect -2035 -964 -1985 -947
rect -2143 -981 -2127 -964
rect -2259 -997 -2127 -981
rect -2001 -981 -1985 -964
rect -1885 -964 -1835 -947
rect -1777 -947 -1577 -900
rect -1777 -964 -1727 -947
rect -1885 -981 -1869 -964
rect -2001 -997 -1869 -981
rect -1743 -981 -1727 -964
rect -1627 -964 -1577 -947
rect -1519 -947 -1319 -900
rect -1519 -964 -1469 -947
rect -1627 -981 -1611 -964
rect -1743 -997 -1611 -981
rect -1485 -981 -1469 -964
rect -1369 -964 -1319 -947
rect -1261 -947 -1061 -900
rect -1261 -964 -1211 -947
rect -1369 -981 -1353 -964
rect -1485 -997 -1353 -981
rect -1227 -981 -1211 -964
rect -1111 -964 -1061 -947
rect -1003 -947 -803 -900
rect -1003 -964 -953 -947
rect -1111 -981 -1095 -964
rect -1227 -997 -1095 -981
rect -969 -981 -953 -964
rect -853 -964 -803 -947
rect -745 -947 -545 -900
rect -745 -964 -695 -947
rect -853 -981 -837 -964
rect -969 -997 -837 -981
rect -711 -981 -695 -964
rect -595 -964 -545 -947
rect -487 -947 -287 -900
rect -487 -964 -437 -947
rect -595 -981 -579 -964
rect -711 -997 -579 -981
rect -453 -981 -437 -964
rect -337 -964 -287 -947
rect -229 -947 -29 -900
rect -229 -964 -179 -947
rect -337 -981 -321 -964
rect -453 -997 -321 -981
rect -195 -981 -179 -964
rect -79 -964 -29 -947
rect 29 -947 229 -900
rect 29 -964 79 -947
rect -79 -981 -63 -964
rect -195 -997 -63 -981
rect 63 -981 79 -964
rect 179 -964 229 -947
rect 287 -947 487 -900
rect 287 -964 337 -947
rect 179 -981 195 -964
rect 63 -997 195 -981
rect 321 -981 337 -964
rect 437 -964 487 -947
rect 545 -947 745 -900
rect 545 -964 595 -947
rect 437 -981 453 -964
rect 321 -997 453 -981
rect 579 -981 595 -964
rect 695 -964 745 -947
rect 803 -947 1003 -900
rect 803 -964 853 -947
rect 695 -981 711 -964
rect 579 -997 711 -981
rect 837 -981 853 -964
rect 953 -964 1003 -947
rect 1061 -947 1261 -900
rect 1061 -964 1111 -947
rect 953 -981 969 -964
rect 837 -997 969 -981
rect 1095 -981 1111 -964
rect 1211 -964 1261 -947
rect 1319 -947 1519 -900
rect 1319 -964 1369 -947
rect 1211 -981 1227 -964
rect 1095 -997 1227 -981
rect 1353 -981 1369 -964
rect 1469 -964 1519 -947
rect 1577 -947 1777 -900
rect 1577 -964 1627 -947
rect 1469 -981 1485 -964
rect 1353 -997 1485 -981
rect 1611 -981 1627 -964
rect 1727 -964 1777 -947
rect 1835 -947 2035 -900
rect 1835 -964 1885 -947
rect 1727 -981 1743 -964
rect 1611 -997 1743 -981
rect 1869 -981 1885 -964
rect 1985 -964 2035 -947
rect 2093 -947 2293 -900
rect 2093 -964 2143 -947
rect 1985 -981 2001 -964
rect 1869 -997 2001 -981
rect 2127 -981 2143 -964
rect 2243 -964 2293 -947
rect 2351 -947 2551 -900
rect 2351 -964 2401 -947
rect 2243 -981 2259 -964
rect 2127 -997 2259 -981
rect 2385 -981 2401 -964
rect 2501 -964 2551 -947
rect 2609 -947 2809 -900
rect 2609 -964 2659 -947
rect 2501 -981 2517 -964
rect 2385 -997 2517 -981
rect 2643 -981 2659 -964
rect 2759 -964 2809 -947
rect 2759 -981 2775 -964
rect 2643 -997 2775 -981
<< polycont >>
rect -2759 947 -2659 981
rect -2501 947 -2401 981
rect -2243 947 -2143 981
rect -1985 947 -1885 981
rect -1727 947 -1627 981
rect -1469 947 -1369 981
rect -1211 947 -1111 981
rect -953 947 -853 981
rect -695 947 -595 981
rect -437 947 -337 981
rect -179 947 -79 981
rect 79 947 179 981
rect 337 947 437 981
rect 595 947 695 981
rect 853 947 953 981
rect 1111 947 1211 981
rect 1369 947 1469 981
rect 1627 947 1727 981
rect 1885 947 1985 981
rect 2143 947 2243 981
rect 2401 947 2501 981
rect 2659 947 2759 981
rect -2759 -981 -2659 -947
rect -2501 -981 -2401 -947
rect -2243 -981 -2143 -947
rect -1985 -981 -1885 -947
rect -1727 -981 -1627 -947
rect -1469 -981 -1369 -947
rect -1211 -981 -1111 -947
rect -953 -981 -853 -947
rect -695 -981 -595 -947
rect -437 -981 -337 -947
rect -179 -981 -79 -947
rect 79 -981 179 -947
rect 337 -981 437 -947
rect 595 -981 695 -947
rect 853 -981 953 -947
rect 1111 -981 1211 -947
rect 1369 -981 1469 -947
rect 1627 -981 1727 -947
rect 1885 -981 1985 -947
rect 2143 -981 2243 -947
rect 2401 -981 2501 -947
rect 2659 -981 2759 -947
<< locali >>
rect -2989 1085 -2893 1119
rect 2893 1085 2989 1119
rect -2989 1023 -2955 1085
rect 2955 1023 2989 1085
rect -2775 947 -2759 981
rect -2659 947 -2643 981
rect -2517 947 -2501 981
rect -2401 947 -2385 981
rect -2259 947 -2243 981
rect -2143 947 -2127 981
rect -2001 947 -1985 981
rect -1885 947 -1869 981
rect -1743 947 -1727 981
rect -1627 947 -1611 981
rect -1485 947 -1469 981
rect -1369 947 -1353 981
rect -1227 947 -1211 981
rect -1111 947 -1095 981
rect -969 947 -953 981
rect -853 947 -837 981
rect -711 947 -695 981
rect -595 947 -579 981
rect -453 947 -437 981
rect -337 947 -321 981
rect -195 947 -179 981
rect -79 947 -63 981
rect 63 947 79 981
rect 179 947 195 981
rect 321 947 337 981
rect 437 947 453 981
rect 579 947 595 981
rect 695 947 711 981
rect 837 947 853 981
rect 953 947 969 981
rect 1095 947 1111 981
rect 1211 947 1227 981
rect 1353 947 1369 981
rect 1469 947 1485 981
rect 1611 947 1627 981
rect 1727 947 1743 981
rect 1869 947 1885 981
rect 1985 947 2001 981
rect 2127 947 2143 981
rect 2243 947 2259 981
rect 2385 947 2401 981
rect 2501 947 2517 981
rect 2643 947 2659 981
rect 2759 947 2775 981
rect -2855 888 -2821 904
rect -2855 -904 -2821 -888
rect -2597 888 -2563 904
rect -2597 -904 -2563 -888
rect -2339 888 -2305 904
rect -2339 -904 -2305 -888
rect -2081 888 -2047 904
rect -2081 -904 -2047 -888
rect -1823 888 -1789 904
rect -1823 -904 -1789 -888
rect -1565 888 -1531 904
rect -1565 -904 -1531 -888
rect -1307 888 -1273 904
rect -1307 -904 -1273 -888
rect -1049 888 -1015 904
rect -1049 -904 -1015 -888
rect -791 888 -757 904
rect -791 -904 -757 -888
rect -533 888 -499 904
rect -533 -904 -499 -888
rect -275 888 -241 904
rect -275 -904 -241 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 241 888 275 904
rect 241 -904 275 -888
rect 499 888 533 904
rect 499 -904 533 -888
rect 757 888 791 904
rect 757 -904 791 -888
rect 1015 888 1049 904
rect 1015 -904 1049 -888
rect 1273 888 1307 904
rect 1273 -904 1307 -888
rect 1531 888 1565 904
rect 1531 -904 1565 -888
rect 1789 888 1823 904
rect 1789 -904 1823 -888
rect 2047 888 2081 904
rect 2047 -904 2081 -888
rect 2305 888 2339 904
rect 2305 -904 2339 -888
rect 2563 888 2597 904
rect 2563 -904 2597 -888
rect 2821 888 2855 904
rect 2821 -904 2855 -888
rect -2775 -981 -2759 -947
rect -2659 -981 -2643 -947
rect -2517 -981 -2501 -947
rect -2401 -981 -2385 -947
rect -2259 -981 -2243 -947
rect -2143 -981 -2127 -947
rect -2001 -981 -1985 -947
rect -1885 -981 -1869 -947
rect -1743 -981 -1727 -947
rect -1627 -981 -1611 -947
rect -1485 -981 -1469 -947
rect -1369 -981 -1353 -947
rect -1227 -981 -1211 -947
rect -1111 -981 -1095 -947
rect -969 -981 -953 -947
rect -853 -981 -837 -947
rect -711 -981 -695 -947
rect -595 -981 -579 -947
rect -453 -981 -437 -947
rect -337 -981 -321 -947
rect -195 -981 -179 -947
rect -79 -981 -63 -947
rect 63 -981 79 -947
rect 179 -981 195 -947
rect 321 -981 337 -947
rect 437 -981 453 -947
rect 579 -981 595 -947
rect 695 -981 711 -947
rect 837 -981 853 -947
rect 953 -981 969 -947
rect 1095 -981 1111 -947
rect 1211 -981 1227 -947
rect 1353 -981 1369 -947
rect 1469 -981 1485 -947
rect 1611 -981 1627 -947
rect 1727 -981 1743 -947
rect 1869 -981 1885 -947
rect 1985 -981 2001 -947
rect 2127 -981 2143 -947
rect 2243 -981 2259 -947
rect 2385 -981 2401 -947
rect 2501 -981 2517 -947
rect 2643 -981 2659 -947
rect 2759 -981 2775 -947
rect -2989 -1085 -2955 -1023
rect 2955 -1085 2989 -1023
rect -2989 -1119 -2893 -1085
rect 2893 -1119 2989 -1085
<< viali >>
rect -2759 947 -2659 981
rect -2501 947 -2401 981
rect -2243 947 -2143 981
rect -1985 947 -1885 981
rect -1727 947 -1627 981
rect -1469 947 -1369 981
rect -1211 947 -1111 981
rect -953 947 -853 981
rect -695 947 -595 981
rect -437 947 -337 981
rect -179 947 -79 981
rect 79 947 179 981
rect 337 947 437 981
rect 595 947 695 981
rect 853 947 953 981
rect 1111 947 1211 981
rect 1369 947 1469 981
rect 1627 947 1727 981
rect 1885 947 1985 981
rect 2143 947 2243 981
rect 2401 947 2501 981
rect 2659 947 2759 981
rect -2855 -888 -2821 888
rect -2597 -888 -2563 888
rect -2339 -888 -2305 888
rect -2081 -888 -2047 888
rect -1823 -888 -1789 888
rect -1565 -888 -1531 888
rect -1307 -888 -1273 888
rect -1049 -888 -1015 888
rect -791 -888 -757 888
rect -533 -888 -499 888
rect -275 -888 -241 888
rect -17 -888 17 888
rect 241 -888 275 888
rect 499 -888 533 888
rect 757 -888 791 888
rect 1015 -888 1049 888
rect 1273 -888 1307 888
rect 1531 -888 1565 888
rect 1789 -888 1823 888
rect 2047 -888 2081 888
rect 2305 -888 2339 888
rect 2563 -888 2597 888
rect 2821 -888 2855 888
rect -2759 -981 -2659 -947
rect -2501 -981 -2401 -947
rect -2243 -981 -2143 -947
rect -1985 -981 -1885 -947
rect -1727 -981 -1627 -947
rect -1469 -981 -1369 -947
rect -1211 -981 -1111 -947
rect -953 -981 -853 -947
rect -695 -981 -595 -947
rect -437 -981 -337 -947
rect -179 -981 -79 -947
rect 79 -981 179 -947
rect 337 -981 437 -947
rect 595 -981 695 -947
rect 853 -981 953 -947
rect 1111 -981 1211 -947
rect 1369 -981 1469 -947
rect 1627 -981 1727 -947
rect 1885 -981 1985 -947
rect 2143 -981 2243 -947
rect 2401 -981 2501 -947
rect 2659 -981 2759 -947
<< metal1 >>
rect -2771 981 -2647 987
rect -2771 947 -2759 981
rect -2659 947 -2647 981
rect -2771 941 -2647 947
rect -2513 981 -2389 987
rect -2513 947 -2501 981
rect -2401 947 -2389 981
rect -2513 941 -2389 947
rect -2255 981 -2131 987
rect -2255 947 -2243 981
rect -2143 947 -2131 981
rect -2255 941 -2131 947
rect -1997 981 -1873 987
rect -1997 947 -1985 981
rect -1885 947 -1873 981
rect -1997 941 -1873 947
rect -1739 981 -1615 987
rect -1739 947 -1727 981
rect -1627 947 -1615 981
rect -1739 941 -1615 947
rect -1481 981 -1357 987
rect -1481 947 -1469 981
rect -1369 947 -1357 981
rect -1481 941 -1357 947
rect -1223 981 -1099 987
rect -1223 947 -1211 981
rect -1111 947 -1099 981
rect -1223 941 -1099 947
rect -965 981 -841 987
rect -965 947 -953 981
rect -853 947 -841 981
rect -965 941 -841 947
rect -707 981 -583 987
rect -707 947 -695 981
rect -595 947 -583 981
rect -707 941 -583 947
rect -449 981 -325 987
rect -449 947 -437 981
rect -337 947 -325 981
rect -449 941 -325 947
rect -191 981 -67 987
rect -191 947 -179 981
rect -79 947 -67 981
rect -191 941 -67 947
rect 67 981 191 987
rect 67 947 79 981
rect 179 947 191 981
rect 67 941 191 947
rect 325 981 449 987
rect 325 947 337 981
rect 437 947 449 981
rect 325 941 449 947
rect 583 981 707 987
rect 583 947 595 981
rect 695 947 707 981
rect 583 941 707 947
rect 841 981 965 987
rect 841 947 853 981
rect 953 947 965 981
rect 841 941 965 947
rect 1099 981 1223 987
rect 1099 947 1111 981
rect 1211 947 1223 981
rect 1099 941 1223 947
rect 1357 981 1481 987
rect 1357 947 1369 981
rect 1469 947 1481 981
rect 1357 941 1481 947
rect 1615 981 1739 987
rect 1615 947 1627 981
rect 1727 947 1739 981
rect 1615 941 1739 947
rect 1873 981 1997 987
rect 1873 947 1885 981
rect 1985 947 1997 981
rect 1873 941 1997 947
rect 2131 981 2255 987
rect 2131 947 2143 981
rect 2243 947 2255 981
rect 2131 941 2255 947
rect 2389 981 2513 987
rect 2389 947 2401 981
rect 2501 947 2513 981
rect 2389 941 2513 947
rect 2647 981 2771 987
rect 2647 947 2659 981
rect 2759 947 2771 981
rect 2647 941 2771 947
rect -2861 888 -2815 900
rect -2861 -888 -2855 888
rect -2821 -888 -2815 888
rect -2861 -900 -2815 -888
rect -2603 888 -2557 900
rect -2603 -888 -2597 888
rect -2563 -888 -2557 888
rect -2603 -900 -2557 -888
rect -2345 888 -2299 900
rect -2345 -888 -2339 888
rect -2305 -888 -2299 888
rect -2345 -900 -2299 -888
rect -2087 888 -2041 900
rect -2087 -888 -2081 888
rect -2047 -888 -2041 888
rect -2087 -900 -2041 -888
rect -1829 888 -1783 900
rect -1829 -888 -1823 888
rect -1789 -888 -1783 888
rect -1829 -900 -1783 -888
rect -1571 888 -1525 900
rect -1571 -888 -1565 888
rect -1531 -888 -1525 888
rect -1571 -900 -1525 -888
rect -1313 888 -1267 900
rect -1313 -888 -1307 888
rect -1273 -888 -1267 888
rect -1313 -900 -1267 -888
rect -1055 888 -1009 900
rect -1055 -888 -1049 888
rect -1015 -888 -1009 888
rect -1055 -900 -1009 -888
rect -797 888 -751 900
rect -797 -888 -791 888
rect -757 -888 -751 888
rect -797 -900 -751 -888
rect -539 888 -493 900
rect -539 -888 -533 888
rect -499 -888 -493 888
rect -539 -900 -493 -888
rect -281 888 -235 900
rect -281 -888 -275 888
rect -241 -888 -235 888
rect -281 -900 -235 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 235 888 281 900
rect 235 -888 241 888
rect 275 -888 281 888
rect 235 -900 281 -888
rect 493 888 539 900
rect 493 -888 499 888
rect 533 -888 539 888
rect 493 -900 539 -888
rect 751 888 797 900
rect 751 -888 757 888
rect 791 -888 797 888
rect 751 -900 797 -888
rect 1009 888 1055 900
rect 1009 -888 1015 888
rect 1049 -888 1055 888
rect 1009 -900 1055 -888
rect 1267 888 1313 900
rect 1267 -888 1273 888
rect 1307 -888 1313 888
rect 1267 -900 1313 -888
rect 1525 888 1571 900
rect 1525 -888 1531 888
rect 1565 -888 1571 888
rect 1525 -900 1571 -888
rect 1783 888 1829 900
rect 1783 -888 1789 888
rect 1823 -888 1829 888
rect 1783 -900 1829 -888
rect 2041 888 2087 900
rect 2041 -888 2047 888
rect 2081 -888 2087 888
rect 2041 -900 2087 -888
rect 2299 888 2345 900
rect 2299 -888 2305 888
rect 2339 -888 2345 888
rect 2299 -900 2345 -888
rect 2557 888 2603 900
rect 2557 -888 2563 888
rect 2597 -888 2603 888
rect 2557 -900 2603 -888
rect 2815 888 2861 900
rect 2815 -888 2821 888
rect 2855 -888 2861 888
rect 2815 -900 2861 -888
rect -2771 -947 -2647 -941
rect -2771 -981 -2759 -947
rect -2659 -981 -2647 -947
rect -2771 -987 -2647 -981
rect -2513 -947 -2389 -941
rect -2513 -981 -2501 -947
rect -2401 -981 -2389 -947
rect -2513 -987 -2389 -981
rect -2255 -947 -2131 -941
rect -2255 -981 -2243 -947
rect -2143 -981 -2131 -947
rect -2255 -987 -2131 -981
rect -1997 -947 -1873 -941
rect -1997 -981 -1985 -947
rect -1885 -981 -1873 -947
rect -1997 -987 -1873 -981
rect -1739 -947 -1615 -941
rect -1739 -981 -1727 -947
rect -1627 -981 -1615 -947
rect -1739 -987 -1615 -981
rect -1481 -947 -1357 -941
rect -1481 -981 -1469 -947
rect -1369 -981 -1357 -947
rect -1481 -987 -1357 -981
rect -1223 -947 -1099 -941
rect -1223 -981 -1211 -947
rect -1111 -981 -1099 -947
rect -1223 -987 -1099 -981
rect -965 -947 -841 -941
rect -965 -981 -953 -947
rect -853 -981 -841 -947
rect -965 -987 -841 -981
rect -707 -947 -583 -941
rect -707 -981 -695 -947
rect -595 -981 -583 -947
rect -707 -987 -583 -981
rect -449 -947 -325 -941
rect -449 -981 -437 -947
rect -337 -981 -325 -947
rect -449 -987 -325 -981
rect -191 -947 -67 -941
rect -191 -981 -179 -947
rect -79 -981 -67 -947
rect -191 -987 -67 -981
rect 67 -947 191 -941
rect 67 -981 79 -947
rect 179 -981 191 -947
rect 67 -987 191 -981
rect 325 -947 449 -941
rect 325 -981 337 -947
rect 437 -981 449 -947
rect 325 -987 449 -981
rect 583 -947 707 -941
rect 583 -981 595 -947
rect 695 -981 707 -947
rect 583 -987 707 -981
rect 841 -947 965 -941
rect 841 -981 853 -947
rect 953 -981 965 -947
rect 841 -987 965 -981
rect 1099 -947 1223 -941
rect 1099 -981 1111 -947
rect 1211 -981 1223 -947
rect 1099 -987 1223 -981
rect 1357 -947 1481 -941
rect 1357 -981 1369 -947
rect 1469 -981 1481 -947
rect 1357 -987 1481 -981
rect 1615 -947 1739 -941
rect 1615 -981 1627 -947
rect 1727 -981 1739 -947
rect 1615 -987 1739 -981
rect 1873 -947 1997 -941
rect 1873 -981 1885 -947
rect 1985 -981 1997 -947
rect 1873 -987 1997 -981
rect 2131 -947 2255 -941
rect 2131 -981 2143 -947
rect 2243 -981 2255 -947
rect 2131 -987 2255 -981
rect 2389 -947 2513 -941
rect 2389 -981 2401 -947
rect 2501 -981 2513 -947
rect 2389 -987 2513 -981
rect 2647 -947 2771 -941
rect 2647 -981 2659 -947
rect 2759 -981 2771 -947
rect 2647 -987 2771 -981
<< properties >>
string FIXED_BBOX -2972 -1102 2972 1102
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 9 l 1 m 1 nf 22 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

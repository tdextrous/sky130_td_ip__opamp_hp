* NGSPICE file created from sky130_td_ip__opamp_hp.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_W75H7K a_n4673_n1200# a_4873_n1200# a_2093_n1264#
+ a_n4099_n1264# w_n5131_n1497# a_4099_n1200# a_745_n1200# a_1577_n1264# a_803_n1264#
+ a_n745_n1264# a_n1003_n1264# a_n545_n1200# a_4157_n1264# a_n3583_n1264# a_3583_n1200#
+ a_1003_n1200# a_n3383_n1200# a_n2867_n1200# a_3641_n1264# a_n2293_n1264# a_2293_n1200#
+ a_n1577_n1200# a_n2093_n1200# a_n4931_n1200# a_2351_n1264# a_n1777_n1264# a_n4357_n1264#
+ a_1777_n1200# a_n29_n1200# a_n4157_n1200# a_1835_n1264# a_4357_n1200# a_n803_n1200#
+ a_4415_n1264# a_n3841_n1264# a_229_n1200# a_n3641_n1200# a_n229_n1264# a_3841_n1200#
+ a_1061_n1264# a_n3067_n1264# a_3067_n1200# a_3125_n1264# a_n2551_n1264# a_n2351_n1200#
+ a_2609_n1264# a_2551_n1200# a_n1835_n1200# a_n4615_n1264# a_4615_n1200# a_n4415_n1200#
+ a_1319_n1264# a_n1261_n1264# a_1261_n1200# a_n1061_n1200# a_3899_n1264# a_287_n1264#
+ a_n3325_n1264# a_n3125_n1200# a_n2809_n1264# a_3325_n1200# a_n2609_n1200# a_2809_n1200#
+ a_n2035_n1264# a_2035_n1200# a_n1519_n1264# a_1519_n1200# a_n1319_n1200# a_487_n1200#
+ a_n3899_n1200# a_4673_n1264# a_545_n1264# a_29_n1264# a_n487_n1264# a_n287_n1200#
+ a_3383_n1264# a_2867_n1264# a_n4873_n1264#
X0 a_3067_n1200# a_2867_n1264# a_2809_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X1 a_1777_n1200# a_1577_n1264# a_1519_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X2 a_2809_n1200# a_2609_n1264# a_2551_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X3 a_n4157_n1200# a_n4357_n1264# a_n4415_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X4 a_1519_n1200# a_1319_n1264# a_1261_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X5 a_4873_n1200# a_4673_n1264# a_4615_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=1.74 ps=12.29 w=12 l=1
X6 a_3583_n1200# a_3383_n1264# a_3325_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X7 a_4615_n1200# a_4415_n1264# a_4357_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X8 a_n2867_n1200# a_n3067_n1264# a_n3125_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X9 a_487_n1200# a_287_n1264# a_229_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X10 a_2293_n1200# a_2093_n1264# a_2035_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X11 a_3325_n1200# a_3125_n1264# a_3067_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X12 a_n287_n1200# a_n487_n1264# a_n545_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X13 a_n2609_n1200# a_n2809_n1264# a_n2867_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X14 a_n1577_n1200# a_n1777_n1264# a_n1835_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X15 a_n29_n1200# a_n229_n1264# a_n287_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X16 a_n4673_n1200# a_n4873_n1264# a_n4931_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=3.48 ps=24.58 w=12 l=1
X17 a_n1319_n1200# a_n1519_n1264# a_n1577_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X18 a_2035_n1200# a_1835_n1264# a_1777_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X19 a_n4415_n1200# a_n4615_n1264# a_n4673_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X20 a_n3383_n1200# a_n3583_n1264# a_n3641_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X21 a_n3125_n1200# a_n3325_n1264# a_n3383_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X22 a_3841_n1200# a_3641_n1264# a_3583_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X23 a_n2093_n1200# a_n2293_n1264# a_n2351_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X24 a_745_n1200# a_545_n1264# a_487_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X25 a_2551_n1200# a_2351_n1264# a_2293_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X26 a_n1835_n1200# a_n2035_n1264# a_n2093_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X27 a_1261_n1200# a_1061_n1264# a_1003_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X28 a_n545_n1200# a_n745_n1264# a_n803_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X29 a_229_n1200# a_29_n1264# a_n29_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X30 a_4099_n1200# a_3899_n1264# a_3841_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X31 a_n3641_n1200# a_n3841_n1264# a_n3899_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X32 a_n2351_n1200# a_n2551_n1264# a_n2609_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X33 a_1003_n1200# a_803_n1264# a_745_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X34 a_n3899_n1200# a_n4099_n1264# a_n4157_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X35 a_n1061_n1200# a_n1261_n1264# a_n1319_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X36 a_4357_n1200# a_4157_n1264# a_4099_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X37 a_n803_n1200# a_n1003_n1264# a_n1061_n1200# w_n5131_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
C0 w_n5131_n1497# a_n2551_n1264# 0.307639f
C1 a_3841_n1200# a_4099_n1200# 0.655843f
C2 a_1061_n1264# w_n5131_n1497# 0.307639f
C3 a_229_n1200# a_487_n1200# 0.655843f
C4 a_n2351_n1200# a_n2551_n1264# 0.26189f
C5 a_545_n1264# w_n5131_n1497# 0.307639f
C6 a_n2093_n1200# a_n1835_n1200# 0.655843f
C7 a_n2093_n1200# a_n2293_n1264# 0.26189f
C8 a_2809_n1200# a_3067_n1200# 0.655843f
C9 w_n5131_n1497# a_1835_n1264# 0.307639f
C10 a_n2035_n1264# a_n2093_n1200# 0.26189f
C11 a_229_n1200# a_n29_n1200# 0.655843f
C12 w_n5131_n1497# a_4873_n1200# 0.69819f
C13 a_3841_n1200# a_3899_n1264# 0.26189f
C14 a_n3125_n1200# a_n2867_n1200# 0.655843f
C15 w_n5131_n1497# a_4157_n1264# 0.307639f
C16 a_n3383_n1200# a_n3325_n1264# 0.26189f
C17 a_n287_n1200# a_n487_n1264# 0.26189f
C18 a_n1261_n1264# w_n5131_n1497# 0.307639f
C19 a_n4873_n1264# a_n4931_n1200# 0.26189f
C20 a_3067_n1200# a_3325_n1200# 0.655843f
C21 a_n1519_n1264# a_n1319_n1200# 0.26189f
C22 a_803_n1264# a_1003_n1200# 0.26189f
C23 a_n3899_n1200# a_n4099_n1264# 0.26189f
C24 a_n3899_n1200# a_n3641_n1200# 0.655843f
C25 a_n2867_n1200# a_n2609_n1200# 0.655843f
C26 w_n5131_n1497# a_n745_n1264# 0.307639f
C27 a_n29_n1200# a_n229_n1264# 0.26189f
C28 a_2293_n1200# a_2351_n1264# 0.26189f
C29 a_3325_n1200# a_3583_n1200# 0.655843f
C30 a_n4157_n1200# a_n4415_n1200# 0.655843f
C31 a_4673_n1264# a_4873_n1200# 0.26189f
C32 a_n4615_n1264# w_n5131_n1497# 0.307639f
C33 w_n5131_n1497# a_n4357_n1264# 0.307639f
C34 w_n5131_n1497# a_n2293_n1264# 0.307639f
C35 a_n1835_n1200# a_n1577_n1200# 0.655843f
C36 a_n2351_n1200# a_n2293_n1264# 0.26189f
C37 a_n2609_n1200# a_n2351_n1200# 0.655843f
C38 a_n2035_n1264# w_n5131_n1497# 0.307639f
C39 a_n1777_n1264# a_n1835_n1200# 0.26189f
C40 a_3125_n1264# a_3067_n1200# 0.26189f
C41 a_2551_n1200# a_2609_n1264# 0.26189f
C42 a_3583_n1200# a_3841_n1200# 0.655843f
C43 a_n1061_n1200# a_n1261_n1264# 0.26189f
C44 a_2809_n1200# a_2609_n1264# 0.26189f
C45 a_1777_n1200# a_1577_n1264# 0.26189f
C46 a_545_n1264# a_487_n1200# 0.26189f
C47 a_n1577_n1200# a_n1319_n1200# 0.655843f
C48 a_3899_n1264# a_4099_n1200# 0.26189f
C49 a_3383_n1264# a_3325_n1200# 0.26189f
C50 a_3125_n1264# w_n5131_n1497# 0.307639f
C51 a_n803_n1200# a_n1003_n1264# 0.26189f
C52 a_1061_n1264# a_1003_n1200# 0.26189f
C53 w_n5131_n1497# a_n487_n1264# 0.307639f
C54 a_3067_n1200# a_2867_n1264# 0.26189f
C55 a_n3641_n1200# a_n3383_n1200# 0.655843f
C56 a_2035_n1200# a_1835_n1264# 0.26189f
C57 a_2351_n1264# w_n5131_n1497# 0.307639f
C58 a_n2867_n1200# a_n3067_n1264# 0.26189f
C59 a_4157_n1264# a_4357_n1200# 0.26189f
C60 a_n4931_n1200# w_n5131_n1497# 0.69819f
C61 a_n4673_n1200# a_n4615_n1264# 0.26189f
C62 a_n3383_n1200# a_n3583_n1264# 0.26189f
C63 a_3641_n1264# a_3583_n1200# 0.26189f
C64 a_3641_n1264# w_n5131_n1497# 0.307639f
C65 a_29_n1264# w_n5131_n1497# 0.307639f
C66 w_n5131_n1497# a_n3067_n1264# 0.307639f
C67 a_n545_n1200# a_n745_n1264# 0.26189f
C68 a_1319_n1264# a_1261_n1200# 0.26189f
C69 a_2293_n1200# a_2093_n1264# 0.26189f
C70 a_2867_n1264# w_n5131_n1497# 0.307639f
C71 a_n2609_n1200# a_n2809_n1264# 0.26189f
C72 a_n1061_n1200# a_n1319_n1200# 0.655843f
C73 a_4415_n1264# a_4615_n1200# 0.26189f
C74 a_29_n1264# a_229_n1200# 0.26189f
C75 a_n4873_n1264# w_n5131_n1497# 0.34286f
C76 a_2809_n1200# a_2551_n1200# 0.655843f
C77 a_n2609_n1200# a_n2551_n1264# 0.26189f
C78 a_287_n1264# w_n5131_n1497# 0.307639f
C79 a_n4157_n1200# a_n4099_n1264# 0.26189f
C80 w_n5131_n1497# a_1577_n1264# 0.307639f
C81 a_n3325_n1264# w_n5131_n1497# 0.307639f
C82 a_287_n1264# a_229_n1200# 0.26189f
C83 a_1319_n1264# w_n5131_n1497# 0.307639f
C84 w_n5131_n1497# a_3899_n1264# 0.307639f
C85 a_n4931_n1200# a_n4673_n1200# 0.655843f
C86 a_n545_n1200# a_n487_n1264# 0.26189f
C87 a_n1519_n1264# w_n5131_n1497# 0.307639f
C88 a_n2351_n1200# a_n2093_n1200# 0.655843f
C89 a_n1061_n1200# a_n803_n1200# 0.655843f
C90 w_n5131_n1497# a_2093_n1264# 0.307639f
C91 a_n3841_n1264# w_n5131_n1497# 0.307639f
C92 a_n1519_n1264# a_n1577_n1200# 0.26189f
C93 a_803_n1264# a_745_n1200# 0.26189f
C94 a_n3641_n1200# a_n3841_n1264# 0.26189f
C95 w_n5131_n1497# a_4415_n1264# 0.307639f
C96 a_n4673_n1200# a_n4415_n1200# 0.655843f
C97 w_n5131_n1497# a_n1003_n1264# 0.307639f
C98 a_n287_n1200# a_n229_n1264# 0.26189f
C99 a_n4873_n1264# a_n4673_n1200# 0.26189f
C100 a_n803_n1200# a_n545_n1200# 0.655843f
C101 a_4673_n1264# a_4615_n1200# 0.26189f
C102 a_n1261_n1264# a_n1319_n1200# 0.26189f
C103 a_29_n1264# a_n29_n1200# 0.26189f
C104 a_n2035_n1264# a_n1835_n1200# 0.26189f
C105 a_2551_n1200# a_2351_n1264# 0.26189f
C106 a_1519_n1200# a_1777_n1200# 0.655843f
C107 a_n3383_n1200# a_n3125_n1200# 0.655843f
C108 a_n545_n1200# a_n287_n1200# 0.655843f
C109 a_1519_n1200# a_1577_n1264# 0.26189f
C110 a_287_n1264# a_487_n1200# 0.26189f
C111 a_4099_n1200# a_4357_n1200# 0.655843f
C112 a_487_n1200# a_745_n1200# 0.655843f
C113 w_n5131_n1497# a_n4099_n1264# 0.307639f
C114 a_n1777_n1264# w_n5131_n1497# 0.307639f
C115 a_1319_n1264# a_1519_n1200# 0.26189f
C116 a_n1777_n1264# a_n1577_n1200# 0.26189f
C117 a_3125_n1264# a_3325_n1200# 0.26189f
C118 a_1777_n1200# a_2035_n1200# 0.655843f
C119 a_n287_n1200# a_n29_n1200# 0.655843f
C120 a_n1061_n1200# a_n1003_n1264# 0.26189f
C121 a_1261_n1200# a_1519_n1200# 0.655843f
C122 a_2809_n1200# a_2867_n1264# 0.26189f
C123 a_1777_n1200# a_1835_n1264# 0.26189f
C124 a_545_n1264# a_745_n1200# 0.26189f
C125 a_n3583_n1264# w_n5131_n1497# 0.307639f
C126 a_803_n1264# w_n5131_n1497# 0.307639f
C127 a_n3125_n1200# a_n3067_n1264# 0.26189f
C128 a_4357_n1200# a_4615_n1200# 0.655843f
C129 a_745_n1200# a_1003_n1200# 0.655843f
C130 a_4157_n1264# a_4099_n1200# 0.26189f
C131 a_4673_n1264# w_n5131_n1497# 0.34286f
C132 a_n3641_n1200# a_n3583_n1264# 0.26189f
C133 a_3383_n1264# a_3583_n1200# 0.26189f
C134 a_2035_n1200# a_2293_n1200# 0.655843f
C135 a_3383_n1264# w_n5131_n1497# 0.307639f
C136 a_n4157_n1200# a_n3899_n1200# 0.655843f
C137 a_n803_n1200# a_n745_n1264# 0.26189f
C138 a_1061_n1264# a_1261_n1200# 0.26189f
C139 w_n5131_n1497# a_n229_n1264# 0.307639f
C140 a_2035_n1200# a_2093_n1264# 0.26189f
C141 a_2609_n1264# w_n5131_n1497# 0.307639f
C142 a_n2867_n1200# a_n2809_n1264# 0.26189f
C143 a_4615_n1200# a_4873_n1200# 0.655843f
C144 a_1003_n1200# a_1261_n1200# 0.655843f
C145 a_4415_n1264# a_4357_n1200# 0.26189f
C146 a_n4415_n1200# a_n4615_n1264# 0.26189f
C147 a_n4415_n1200# a_n4357_n1264# 0.26189f
C148 a_3641_n1264# a_3841_n1200# 0.26189f
C149 a_2293_n1200# a_2551_n1200# 0.655843f
C150 a_n3125_n1200# a_n3325_n1264# 0.26189f
C151 w_n5131_n1497# a_n2809_n1264# 0.307639f
C152 a_n4157_n1200# a_n4357_n1264# 0.26189f
C153 a_n3899_n1200# a_n3841_n1264# 0.26189f
C154 a_4873_n1200# 0 0.58762f
C155 a_4615_n1200# 0 0.335348f
C156 a_4357_n1200# 0 0.335348f
C157 a_4099_n1200# 0 0.335348f
C158 a_3841_n1200# 0 0.335348f
C159 a_3583_n1200# 0 0.335348f
C160 a_3325_n1200# 0 0.335348f
C161 a_3067_n1200# 0 0.335348f
C162 a_2809_n1200# 0 0.335348f
C163 a_2551_n1200# 0 0.335348f
C164 a_2293_n1200# 0 0.335348f
C165 a_2035_n1200# 0 0.335348f
C166 a_1777_n1200# 0 0.335348f
C167 a_1519_n1200# 0 0.335348f
C168 a_1261_n1200# 0 0.335348f
C169 a_1003_n1200# 0 0.335348f
C170 a_745_n1200# 0 0.335348f
C171 a_487_n1200# 0 0.335348f
C172 a_229_n1200# 0 0.335348f
C173 a_n29_n1200# 0 0.335348f
C174 a_n287_n1200# 0 0.335348f
C175 a_n545_n1200# 0 0.335348f
C176 a_n803_n1200# 0 0.335348f
C177 a_n1061_n1200# 0 0.335348f
C178 a_n1319_n1200# 0 0.335348f
C179 a_n1577_n1200# 0 0.335348f
C180 a_n1835_n1200# 0 0.335348f
C181 a_n2093_n1200# 0 0.335348f
C182 a_n2351_n1200# 0 0.335348f
C183 a_n2609_n1200# 0 0.335348f
C184 a_n2867_n1200# 0 0.335348f
C185 a_n3125_n1200# 0 0.335348f
C186 a_n3383_n1200# 0 0.335348f
C187 a_n3641_n1200# 0 0.335348f
C188 a_n3899_n1200# 0 0.335348f
C189 a_n4157_n1200# 0 0.335348f
C190 a_n4415_n1200# 0 0.335348f
C191 a_n4673_n1200# 0 0.335348f
C192 a_n4931_n1200# 0 0.58762f
C193 a_4673_n1264# 0 0.253452f
C194 a_4415_n1264# 0 0.231023f
C195 a_4157_n1264# 0 0.231023f
C196 a_3899_n1264# 0 0.231023f
C197 a_3641_n1264# 0 0.231023f
C198 a_3383_n1264# 0 0.231023f
C199 a_3125_n1264# 0 0.231023f
C200 a_2867_n1264# 0 0.231023f
C201 a_2609_n1264# 0 0.231023f
C202 a_2351_n1264# 0 0.231023f
C203 a_2093_n1264# 0 0.231023f
C204 a_1835_n1264# 0 0.231023f
C205 a_1577_n1264# 0 0.231023f
C206 a_1319_n1264# 0 0.231023f
C207 a_1061_n1264# 0 0.231023f
C208 a_803_n1264# 0 0.231023f
C209 a_545_n1264# 0 0.231023f
C210 a_287_n1264# 0 0.231023f
C211 a_29_n1264# 0 0.231023f
C212 a_n229_n1264# 0 0.231023f
C213 a_n487_n1264# 0 0.231023f
C214 a_n745_n1264# 0 0.231023f
C215 a_n1003_n1264# 0 0.231023f
C216 a_n1261_n1264# 0 0.231023f
C217 a_n1519_n1264# 0 0.231023f
C218 a_n1777_n1264# 0 0.231023f
C219 a_n2035_n1264# 0 0.231023f
C220 a_n2293_n1264# 0 0.231023f
C221 a_n2551_n1264# 0 0.231023f
C222 a_n2809_n1264# 0 0.231023f
C223 a_n3067_n1264# 0 0.231023f
C224 a_n3325_n1264# 0 0.231023f
C225 a_n3583_n1264# 0 0.231023f
C226 a_n3841_n1264# 0 0.231023f
C227 a_n4099_n1264# 0 0.231023f
C228 a_n4357_n1264# 0 0.231023f
C229 a_n4615_n1264# 0 0.231023f
C230 a_n4873_n1264# 0 0.253452f
C231 w_n5131_n1497# 0 99.8345f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_CVG6CD a_50_n400# w_n308_n697# a_n50_n464# a_n108_n400#
X0 a_50_n400# a_n50_n464# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
C0 w_n308_n697# a_50_n400# 0.249352f
C1 w_n308_n697# a_n50_n464# 0.259326f
C2 w_n308_n697# a_n108_n400# 0.249352f
C3 a_n108_n400# a_50_n400# 0.357178f
C4 a_50_n400# 0 0.180042f
C5 a_n108_n400# 0 0.180042f
C6 a_n50_n464# 0 0.148749f
C7 w_n308_n697# 0 3.40572f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_WKXP7K a_n4673_n1200# a_4873_n1200# a_4931_n1264#
+ a_2093_n1264# a_n4099_n1264# a_4099_n1200# a_745_n1200# a_1577_n1264# a_803_n1264#
+ a_n745_n1264# a_n1003_n1264# a_n545_n1200# a_4157_n1264# a_n3583_n1264# a_3583_n1200#
+ a_1003_n1200# a_n3383_n1200# a_n2867_n1200# a_3641_n1264# a_n2293_n1264# a_2293_n1200#
+ a_n1577_n1200# a_n2093_n1200# a_n4931_n1200# a_2351_n1264# a_n1777_n1264# a_n4357_n1264#
+ a_1777_n1200# a_n29_n1200# a_n4157_n1200# a_1835_n1264# a_4357_n1200# a_n803_n1200#
+ a_4415_n1264# a_n3841_n1264# a_229_n1200# a_n3641_n1200# a_n229_n1264# a_3841_n1200#
+ a_1061_n1264# a_n3067_n1264# a_3067_n1200# a_3125_n1264# a_n2551_n1264# a_n2351_n1200#
+ a_2609_n1264# a_n5131_n1264# w_n5389_n1497# a_5131_n1200# a_2551_n1200# a_n1835_n1200#
+ a_n4615_n1264# a_4615_n1200# a_n4415_n1200# a_1319_n1264# a_n1261_n1264# a_1261_n1200#
+ a_n1061_n1200# a_3899_n1264# a_287_n1264# a_n3325_n1264# a_n3125_n1200# a_n2809_n1264#
+ a_3325_n1200# a_n2609_n1200# a_2809_n1200# a_n2035_n1264# a_2035_n1200# a_n1519_n1264#
+ a_1519_n1200# a_n1319_n1200# a_487_n1200# a_n3899_n1200# a_4673_n1264# a_545_n1264#
+ a_29_n1264# a_n487_n1264# a_n287_n1200# a_3383_n1264# a_n5189_n1200# a_2867_n1264#
+ a_n4873_n1264#
X0 a_3067_n1200# a_2867_n1264# a_2809_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X1 a_1777_n1200# a_1577_n1264# a_1519_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X2 a_2809_n1200# a_2609_n1264# a_2551_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X3 a_n4157_n1200# a_n4357_n1264# a_n4415_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X4 a_1519_n1200# a_1319_n1264# a_1261_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X5 a_4873_n1200# a_4673_n1264# a_4615_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X6 a_3583_n1200# a_3383_n1264# a_3325_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X7 a_4615_n1200# a_4415_n1264# a_4357_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X8 a_n2867_n1200# a_n3067_n1264# a_n3125_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X9 a_487_n1200# a_287_n1264# a_229_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X10 a_2293_n1200# a_2093_n1264# a_2035_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X11 a_3325_n1200# a_3125_n1264# a_3067_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X12 a_n287_n1200# a_n487_n1264# a_n545_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X13 a_n2609_n1200# a_n2809_n1264# a_n2867_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X14 a_n1577_n1200# a_n1777_n1264# a_n1835_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X15 a_n29_n1200# a_n229_n1264# a_n287_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X16 a_n4673_n1200# a_n4873_n1264# a_n4931_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X17 a_n1319_n1200# a_n1519_n1264# a_n1577_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X18 a_2035_n1200# a_1835_n1264# a_1777_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X19 a_5131_n1200# a_4931_n1264# a_4873_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=1.74 ps=12.29 w=12 l=1
X20 a_n4415_n1200# a_n4615_n1264# a_n4673_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X21 a_n3383_n1200# a_n3583_n1264# a_n3641_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X22 a_n3125_n1200# a_n3325_n1264# a_n3383_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X23 a_3841_n1200# a_3641_n1264# a_3583_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X24 a_n2093_n1200# a_n2293_n1264# a_n2351_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X25 a_745_n1200# a_545_n1264# a_487_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X26 a_2551_n1200# a_2351_n1264# a_2293_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X27 a_n1835_n1200# a_n2035_n1264# a_n2093_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X28 a_n4931_n1200# a_n5131_n1264# a_n5189_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=3.48 ps=24.58 w=12 l=1
X29 a_1261_n1200# a_1061_n1264# a_1003_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X30 a_n545_n1200# a_n745_n1264# a_n803_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X31 a_229_n1200# a_29_n1264# a_n29_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X32 a_4099_n1200# a_3899_n1264# a_3841_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X33 a_n3641_n1200# a_n3841_n1264# a_n3899_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X34 a_n2351_n1200# a_n2551_n1264# a_n2609_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X35 a_1003_n1200# a_803_n1264# a_745_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X36 a_n3899_n1200# a_n4099_n1264# a_n4157_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X37 a_n1061_n1200# a_n1261_n1264# a_n1319_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X38 a_4357_n1200# a_4157_n1264# a_4099_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
X39 a_n803_n1200# a_n1003_n1264# a_n1061_n1200# w_n5389_n1497# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.29 as=1.74 ps=12.29 w=12 l=1
C0 a_n4157_n1200# a_n3899_n1200# 0.655843f
C1 a_n545_n1200# a_n287_n1200# 0.655843f
C2 w_n5389_n1497# a_n4615_n1264# 0.307639f
C3 a_n3899_n1200# a_n4099_n1264# 0.26189f
C4 a_n1577_n1200# a_n1319_n1200# 0.655843f
C5 a_1777_n1200# a_1835_n1264# 0.26189f
C6 a_n2293_n1264# a_n2093_n1200# 0.26189f
C7 a_2551_n1200# a_2609_n1264# 0.26189f
C8 a_n487_n1264# a_n287_n1200# 0.26189f
C9 a_n3841_n1264# a_n3899_n1200# 0.26189f
C10 w_n5389_n1497# a_n4099_n1264# 0.307639f
C11 a_n1835_n1200# a_n1777_n1264# 0.26189f
C12 a_n1519_n1264# a_n1577_n1200# 0.26189f
C13 a_3067_n1200# a_2867_n1264# 0.26189f
C14 a_n2035_n1264# a_n2093_n1200# 0.26189f
C15 a_1519_n1200# a_1319_n1264# 0.26189f
C16 a_n4673_n1200# a_n4873_n1264# 0.26189f
C17 a_n3841_n1264# w_n5389_n1497# 0.307639f
C18 a_n29_n1200# a_29_n1264# 0.26189f
C19 a_n2809_n1264# w_n5389_n1497# 0.307639f
C20 w_n5389_n1497# a_1577_n1264# 0.307639f
C21 a_229_n1200# a_29_n1264# 0.26189f
C22 a_3325_n1200# a_3383_n1264# 0.26189f
C23 a_n29_n1200# a_n287_n1200# 0.655843f
C24 a_n29_n1200# a_n229_n1264# 0.26189f
C25 a_745_n1200# a_803_n1264# 0.26189f
C26 w_n5389_n1497# a_3383_n1264# 0.307639f
C27 w_n5389_n1497# a_2867_n1264# 0.307639f
C28 w_n5389_n1497# a_4415_n1264# 0.307639f
C29 a_3841_n1200# a_4099_n1200# 0.655843f
C30 a_3899_n1264# w_n5389_n1497# 0.307639f
C31 a_3899_n1264# a_3841_n1200# 0.26189f
C32 a_n2609_n1200# a_n2351_n1200# 0.655843f
C33 a_n2867_n1200# a_n2809_n1264# 0.26189f
C34 w_n5389_n1497# a_n487_n1264# 0.307639f
C35 a_n1003_n1264# a_n1061_n1200# 0.26189f
C36 a_n1061_n1200# a_n1319_n1200# 0.655843f
C37 a_745_n1200# a_487_n1200# 0.655843f
C38 a_n2551_n1264# a_n2351_n1200# 0.26189f
C39 a_4357_n1200# a_4415_n1264# 0.26189f
C40 a_4357_n1200# a_4099_n1200# 0.655843f
C41 a_n3583_n1264# a_n3383_n1200# 0.26189f
C42 w_n5389_n1497# a_n5131_n1264# 0.34286f
C43 a_n5189_n1200# a_n4931_n1200# 0.655843f
C44 a_2551_n1200# a_2293_n1200# 0.655843f
C45 a_2809_n1200# a_2867_n1264# 0.26189f
C46 a_4615_n1200# a_4415_n1264# 0.26189f
C47 a_487_n1200# a_287_n1264# 0.26189f
C48 a_n3583_n1264# w_n5389_n1497# 0.307639f
C49 a_229_n1200# a_487_n1200# 0.655843f
C50 w_n5389_n1497# a_4157_n1264# 0.307639f
C51 a_n545_n1200# a_n803_n1200# 0.655843f
C52 w_n5389_n1497# a_287_n1264# 0.307639f
C53 w_n5389_n1497# a_n1777_n1264# 0.307639f
C54 a_n3841_n1264# a_n3641_n1200# 0.26189f
C55 a_2809_n1200# a_2551_n1200# 0.655843f
C56 a_n2609_n1200# a_n2551_n1264# 0.26189f
C57 a_n5189_n1200# a_n5131_n1264# 0.26189f
C58 a_n4415_n1200# a_n4615_n1264# 0.26189f
C59 a_545_n1264# a_487_n1200# 0.26189f
C60 a_n1519_n1264# a_n1319_n1200# 0.26189f
C61 a_1319_n1264# a_1261_n1200# 0.26189f
C62 a_4357_n1200# a_4157_n1264# 0.26189f
C63 a_1777_n1200# a_2035_n1200# 0.655843f
C64 a_545_n1264# w_n5389_n1497# 0.307639f
C65 a_n287_n1200# a_n229_n1264# 0.26189f
C66 a_3325_n1200# a_3583_n1200# 0.655843f
C67 w_n5389_n1497# a_n745_n1264# 0.307639f
C68 a_1519_n1200# a_1577_n1264# 0.26189f
C69 a_n4157_n1200# a_n4099_n1264# 0.26189f
C70 a_n4415_n1200# a_n4157_n1200# 0.655843f
C71 a_2551_n1200# a_2351_n1264# 0.26189f
C72 a_1261_n1200# a_1003_n1200# 0.655843f
C73 a_745_n1200# a_1003_n1200# 0.655843f
C74 w_n5389_n1497# a_1061_n1264# 0.307639f
C75 a_2093_n1264# a_2293_n1200# 0.26189f
C76 a_2093_n1264# w_n5389_n1497# 0.307639f
C77 a_3841_n1200# a_3583_n1200# 0.655843f
C78 w_n5389_n1497# a_1835_n1264# 0.307639f
C79 w_n5389_n1497# a_n4873_n1264# 0.307639f
C80 w_n5389_n1497# a_2609_n1264# 0.307639f
C81 a_n3325_n1264# a_n3383_n1200# 0.26189f
C82 w_n5389_n1497# a_29_n1264# 0.307639f
C83 a_n1003_n1264# w_n5389_n1497# 0.307639f
C84 a_n1061_n1200# a_n1261_n1264# 0.26189f
C85 a_2093_n1264# a_2035_n1200# 0.26189f
C86 a_1519_n1200# a_1261_n1200# 0.655843f
C87 w_n5389_n1497# a_n4357_n1264# 0.307639f
C88 w_n5389_n1497# a_5131_n1200# 0.69819f
C89 a_n3583_n1264# a_n3641_n1200# 0.26189f
C90 w_n5389_n1497# a_n3325_n1264# 0.307639f
C91 w_n5389_n1497# a_n2551_n1264# 0.307639f
C92 a_4931_n1264# a_5131_n1200# 0.26189f
C93 a_n2093_n1200# a_n2351_n1200# 0.655843f
C94 a_1519_n1200# a_1777_n1200# 0.655843f
C95 a_1835_n1264# a_2035_n1200# 0.26189f
C96 a_n2293_n1264# a_n2351_n1200# 0.26189f
C97 a_n803_n1200# a_n745_n1264# 0.26189f
C98 w_n5389_n1497# a_n229_n1264# 0.307639f
C99 a_2809_n1200# a_2609_n1264# 0.26189f
C100 a_1061_n1264# a_1003_n1200# 0.26189f
C101 a_n1519_n1264# w_n5389_n1497# 0.307639f
C102 a_3067_n1200# a_3325_n1200# 0.655843f
C103 a_n1061_n1200# a_n803_n1200# 0.655843f
C104 a_n1835_n1200# a_n2093_n1200# 0.655843f
C105 a_n2867_n1200# a_n2609_n1200# 0.655843f
C106 a_n1261_n1264# a_n1319_n1200# 0.26189f
C107 a_4673_n1264# w_n5389_n1497# 0.307639f
C108 a_n3125_n1200# a_n3325_n1264# 0.26189f
C109 w_n5389_n1497# a_803_n1264# 0.307639f
C110 a_n4673_n1200# a_n4615_n1264# 0.26189f
C111 a_3583_n1200# a_3641_n1264# 0.26189f
C112 a_3899_n1264# a_4099_n1200# 0.26189f
C113 a_n545_n1200# a_n487_n1264# 0.26189f
C114 a_3125_n1264# a_3067_n1200# 0.26189f
C115 a_n1835_n1200# a_n2035_n1264# 0.26189f
C116 a_n1003_n1264# a_n803_n1200# 0.26189f
C117 a_n5131_n1264# a_n4931_n1200# 0.26189f
C118 a_2809_n1200# a_3067_n1200# 0.655843f
C119 a_1777_n1200# a_1577_n1264# 0.26189f
C120 a_4873_n1200# a_5131_n1200# 0.655843f
C121 a_n4415_n1200# a_n4673_n1200# 0.655843f
C122 a_4615_n1200# a_4673_n1264# 0.26189f
C123 a_4931_n1264# w_n5389_n1497# 0.34286f
C124 a_n3125_n1200# a_n3383_n1200# 0.655843f
C125 a_3125_n1264# a_3325_n1200# 0.26189f
C126 a_3125_n1264# w_n5389_n1497# 0.307639f
C127 a_1003_n1200# a_803_n1264# 0.26189f
C128 a_n4931_n1200# a_n4673_n1200# 0.655843f
C129 w_n5389_n1497# a_n1261_n1264# 0.307639f
C130 a_4673_n1264# a_4873_n1200# 0.26189f
C131 a_4157_n1264# a_4099_n1200# 0.26189f
C132 a_2035_n1200# a_2293_n1200# 0.655843f
C133 a_n5189_n1200# w_n5389_n1497# 0.69819f
C134 a_1319_n1264# w_n5389_n1497# 0.307639f
C135 w_n5389_n1497# a_n3067_n1264# 0.307639f
C136 a_n1577_n1200# a_n1777_n1264# 0.26189f
C137 a_n545_n1200# a_n745_n1264# 0.26189f
C138 a_4615_n1200# a_4357_n1200# 0.655843f
C139 a_2351_n1264# a_2293_n1200# 0.26189f
C140 w_n5389_n1497# a_2351_n1264# 0.307639f
C141 a_n4157_n1200# a_n4357_n1264# 0.26189f
C142 a_n2293_n1264# w_n5389_n1497# 0.307639f
C143 a_n2867_n1200# a_n3125_n1200# 0.655843f
C144 a_n3641_n1200# a_n3383_n1200# 0.655843f
C145 a_n3899_n1200# a_n3641_n1200# 0.655843f
C146 a_n4415_n1200# a_n4357_n1264# 0.26189f
C147 a_n4931_n1200# a_n4873_n1264# 0.26189f
C148 a_3583_n1200# a_3383_n1264# 0.26189f
C149 a_4931_n1264# a_4873_n1200# 0.26189f
C150 a_n3125_n1200# a_n3067_n1264# 0.26189f
C151 a_n2867_n1200# a_n3067_n1264# 0.26189f
C152 w_n5389_n1497# a_3641_n1264# 0.307639f
C153 a_n2809_n1264# a_n2609_n1200# 0.26189f
C154 a_3841_n1200# a_3641_n1264# 0.26189f
C155 a_545_n1264# a_745_n1200# 0.26189f
C156 w_n5389_n1497# a_n2035_n1264# 0.307639f
C157 a_n1835_n1200# a_n1577_n1200# 0.655843f
C158 a_n29_n1200# a_229_n1200# 0.655843f
C159 a_1261_n1200# a_1061_n1264# 0.26189f
C160 a_229_n1200# a_287_n1264# 0.26189f
C161 a_4615_n1200# a_4873_n1200# 0.655843f
C162 a_5131_n1200# 0 0.58762f
C163 a_4873_n1200# 0 0.335348f
C164 a_4615_n1200# 0 0.335348f
C165 a_4357_n1200# 0 0.335348f
C166 a_4099_n1200# 0 0.335348f
C167 a_3841_n1200# 0 0.335348f
C168 a_3583_n1200# 0 0.335348f
C169 a_3325_n1200# 0 0.335348f
C170 a_3067_n1200# 0 0.335348f
C171 a_2809_n1200# 0 0.335348f
C172 a_2551_n1200# 0 0.335348f
C173 a_2293_n1200# 0 0.335348f
C174 a_2035_n1200# 0 0.335348f
C175 a_1777_n1200# 0 0.335348f
C176 a_1519_n1200# 0 0.335348f
C177 a_1261_n1200# 0 0.335348f
C178 a_1003_n1200# 0 0.335348f
C179 a_745_n1200# 0 0.335348f
C180 a_487_n1200# 0 0.335348f
C181 a_229_n1200# 0 0.335348f
C182 a_n29_n1200# 0 0.335348f
C183 a_n287_n1200# 0 0.335348f
C184 a_n545_n1200# 0 0.335348f
C185 a_n803_n1200# 0 0.335348f
C186 a_n1061_n1200# 0 0.335348f
C187 a_n1319_n1200# 0 0.335348f
C188 a_n1577_n1200# 0 0.335348f
C189 a_n1835_n1200# 0 0.335348f
C190 a_n2093_n1200# 0 0.335348f
C191 a_n2351_n1200# 0 0.335348f
C192 a_n2609_n1200# 0 0.335348f
C193 a_n2867_n1200# 0 0.335348f
C194 a_n3125_n1200# 0 0.335348f
C195 a_n3383_n1200# 0 0.335348f
C196 a_n3641_n1200# 0 0.335348f
C197 a_n3899_n1200# 0 0.335348f
C198 a_n4157_n1200# 0 0.335348f
C199 a_n4415_n1200# 0 0.335348f
C200 a_n4673_n1200# 0 0.335348f
C201 a_n4931_n1200# 0 0.335348f
C202 a_n5189_n1200# 0 0.58762f
C203 a_4931_n1264# 0 0.253452f
C204 a_4673_n1264# 0 0.231023f
C205 a_4415_n1264# 0 0.231023f
C206 a_4157_n1264# 0 0.231023f
C207 a_3899_n1264# 0 0.231023f
C208 a_3641_n1264# 0 0.231023f
C209 a_3383_n1264# 0 0.231023f
C210 a_3125_n1264# 0 0.231023f
C211 a_2867_n1264# 0 0.231023f
C212 a_2609_n1264# 0 0.231023f
C213 a_2351_n1264# 0 0.231023f
C214 a_2093_n1264# 0 0.231023f
C215 a_1835_n1264# 0 0.231023f
C216 a_1577_n1264# 0 0.231023f
C217 a_1319_n1264# 0 0.231023f
C218 a_1061_n1264# 0 0.231023f
C219 a_803_n1264# 0 0.231023f
C220 a_545_n1264# 0 0.231023f
C221 a_287_n1264# 0 0.231023f
C222 a_29_n1264# 0 0.231023f
C223 a_n229_n1264# 0 0.231023f
C224 a_n487_n1264# 0 0.231023f
C225 a_n745_n1264# 0 0.231023f
C226 a_n1003_n1264# 0 0.231023f
C227 a_n1261_n1264# 0 0.231023f
C228 a_n1519_n1264# 0 0.231023f
C229 a_n1777_n1264# 0 0.231023f
C230 a_n2035_n1264# 0 0.231023f
C231 a_n2293_n1264# 0 0.231023f
C232 a_n2551_n1264# 0 0.231023f
C233 a_n2809_n1264# 0 0.231023f
C234 a_n3067_n1264# 0 0.231023f
C235 a_n3325_n1264# 0 0.231023f
C236 a_n3583_n1264# 0 0.231023f
C237 a_n3841_n1264# 0 0.231023f
C238 a_n4099_n1264# 0 0.231023f
C239 a_n4357_n1264# 0 0.231023f
C240 a_n4615_n1264# 0 0.231023f
C241 a_n4873_n1264# 0 0.231023f
C242 a_n5131_n1264# 0 0.253452f
C243 w_n5389_n1497# 0 0.10479p
.ends

.subckt sky130_fd_pr__nfet_01v8_6H2JYD a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_15_n100# a_n73_n100# 0.162113f
C1 a_15_n100# a_n175_n274# 0.131704f
C2 a_n73_n100# a_n175_n274# 0.131704f
C3 a_n33_n188# a_n175_n274# 0.34289f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CTEUHA a_50_n200# a_n242_n422# a_n108_n200# a_n50_n288#
X0 a_50_n200# a_n50_n288# a_n108_n200# a_n242_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
C0 a_50_n200# a_n108_n200# 0.17948f
C1 a_50_n200# a_n242_n422# 0.231051f
C2 a_n108_n200# a_n242_n422# 0.231051f
C3 a_n50_n288# a_n242_n422# 0.428135f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_HQ4STX w_n358_n597# a_n158_n300# a_n100_n364#
+ a_100_n300#
X0 a_100_n300# a_n100_n364# a_n158_n300# w_n358_n597# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
C0 w_n358_n597# a_n100_n364# 0.378082f
C1 a_n158_n300# w_n358_n597# 0.193235f
C2 a_100_n300# w_n358_n597# 0.193235f
C3 a_100_n300# a_n158_n300# 0.164742f
C4 a_100_n300# 0 0.153252f
C5 a_n158_n300# 0 0.153252f
C6 a_n100_n364# 0 0.25371f
C7 w_n358_n597# 0 3.35808f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YJ3VXJ a_n287_n255# a_n345_n200# a_345_n255#
+ a_n445_n255# a_129_n200# a_n503_n200# a_287_n200# a_445_n200# a_n637_n422# a_n29_n200#
+ a_29_n255# a_n187_n200# a_n129_n255# a_187_n255#
X0 a_n187_n200# a_n287_n255# a_n345_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X1 a_287_n200# a_187_n255# a_129_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X2 a_n345_n200# a_n445_n255# a_n503_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X3 a_129_n200# a_29_n255# a_n29_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
X4 a_445_n200# a_345_n255# a_287_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X5 a_n29_n200# a_n129_n255# a_n187_n200# a_n637_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.5
C0 a_129_n200# a_287_n200# 0.17948f
C1 a_129_n200# a_n29_n200# 0.17948f
C2 a_n345_n200# a_n503_n200# 0.17948f
C3 a_n345_n200# a_n187_n200# 0.17948f
C4 a_445_n200# a_287_n200# 0.17948f
C5 a_n187_n200# a_n29_n200# 0.17948f
C6 a_445_n200# a_n637_n422# 0.231051f
C7 a_n503_n200# a_n637_n422# 0.231051f
C8 a_345_n255# a_n637_n422# 0.33085f
C9 a_187_n255# a_n637_n422# 0.272102f
C10 a_29_n255# a_n637_n422# 0.272102f
C11 a_n129_n255# a_n637_n422# 0.272102f
C12 a_n287_n255# a_n637_n422# 0.272102f
C13 a_n445_n255# a_n637_n422# 0.33085f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J a_1519_n450# a_n803_n450# a_n2093_n450#
+ a_n2551_n505# a_1261_n450# a_29_n505# a_n1777_n505# a_n3067_n505# a_n1319_n450#
+ a_n287_n450# a_n1061_n450# a_2867_n505# a_n745_n505# a_2809_n450# a_803_n505# a_n2035_n505#
+ a_745_n450# a_n3383_n450# a_2551_n450# a_3125_n505# a_1835_n505# a_3067_n450# a_1777_n450#
+ a_n2609_n450# a_n229_n505# a_n1003_n505# a_n2351_n450# a_287_n505# a_2093_n505#
+ a_229_n450# a_n1577_n450# a_n3325_n505# a_2035_n450# a_1319_n505# a_n545_n450# a_1061_n505#
+ a_n2293_n505# a_n3517_n672# a_1003_n450# a_n1519_n505# a_n2867_n450# a_n487_n505#
+ a_3325_n450# a_n1261_n505# a_2609_n505# a_n29_n450# a_545_n505# a_487_n450# a_2351_n505#
+ a_2293_n450# a_n1835_n450# a_n3125_n450# a_1577_n505# a_n2809_n505#
X0 a_n2351_n450# a_n2551_n505# a_n2609_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X1 a_n2093_n450# a_n2293_n505# a_n2351_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X2 a_229_n450# a_29_n505# a_n29_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X3 a_n29_n450# a_n229_n505# a_n287_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X4 a_3067_n450# a_2867_n505# a_2809_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X5 a_n1319_n450# a_n1519_n505# a_n1577_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X6 a_n545_n450# a_n745_n505# a_n803_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X7 a_2551_n450# a_2351_n505# a_2293_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X8 a_n3125_n450# a_n3325_n505# a_n3383_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=1
X9 a_n287_n450# a_n487_n505# a_n545_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X10 a_2293_n450# a_2093_n505# a_2035_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X11 a_n2867_n450# a_n3067_n505# a_n3125_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X12 a_n803_n450# a_n1003_n505# a_n1061_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X13 a_n1577_n450# a_n1777_n505# a_n1835_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X14 a_1519_n450# a_1319_n505# a_1261_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X15 a_n1061_n450# a_n1261_n505# a_n1319_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X16 a_3325_n450# a_3125_n505# a_3067_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=1
X17 a_1003_n450# a_803_n505# a_745_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X18 a_745_n450# a_545_n505# a_487_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X19 a_487_n450# a_287_n505# a_229_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X20 a_2035_n450# a_1835_n505# a_1777_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X21 a_n2609_n450# a_n2809_n505# a_n2867_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X22 a_1777_n450# a_1577_n505# a_1519_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X23 a_1261_n450# a_1061_n505# a_1003_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X24 a_n1835_n450# a_n2035_n505# a_n2093_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X25 a_2809_n450# a_2609_n505# a_2551_n450# a_n3517_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
C0 a_n487_n505# a_n287_n450# 0.101608f
C1 a_n1777_n505# a_n1835_n450# 0.101608f
C2 a_n229_n505# a_n29_n450# 0.101608f
C3 a_3125_n505# a_3325_n450# 0.101608f
C4 a_n2351_n450# a_n2293_n505# 0.101608f
C5 a_2551_n450# a_2609_n505# 0.101608f
C6 a_n1577_n450# a_n1319_n450# 0.246592f
C7 a_2551_n450# a_2809_n450# 0.246592f
C8 a_2809_n450# a_2609_n505# 0.101608f
C9 a_n2809_n505# a_n2609_n450# 0.101608f
C10 a_1261_n450# a_1519_n450# 0.246592f
C11 a_2551_n450# a_2351_n505# 0.101608f
C12 a_n2867_n450# a_n3125_n450# 0.246592f
C13 a_1577_n505# a_1519_n450# 0.101608f
C14 a_803_n505# a_1003_n450# 0.101608f
C15 a_n1319_n450# a_n1261_n505# 0.101608f
C16 a_3067_n450# a_3325_n450# 0.246592f
C17 a_n803_n450# a_n1061_n450# 0.246592f
C18 a_n1577_n450# a_n1519_n505# 0.101608f
C19 a_n2093_n450# a_n2035_n505# 0.101608f
C20 a_2867_n505# a_3067_n450# 0.101608f
C21 a_n3125_n450# a_n3383_n450# 0.246592f
C22 a_29_n505# a_n29_n450# 0.101608f
C23 a_229_n450# a_287_n505# 0.101608f
C24 a_n1319_n450# a_n1519_n505# 0.101608f
C25 a_545_n505# a_487_n450# 0.101608f
C26 a_2551_n450# a_2293_n450# 0.246592f
C27 a_29_n505# a_229_n450# 0.101608f
C28 a_n1777_n505# a_n1577_n450# 0.101608f
C29 a_n287_n450# a_n229_n505# 0.101608f
C30 a_n745_n505# a_n803_n450# 0.101608f
C31 a_2293_n450# a_2351_n505# 0.101608f
C32 a_n1003_n505# a_n1061_n450# 0.101608f
C33 a_n3125_n450# a_n3325_n505# 0.101608f
C34 a_229_n450# a_n29_n450# 0.246592f
C35 a_3067_n450# a_2809_n450# 0.246592f
C36 a_287_n505# a_487_n450# 0.101608f
C37 a_n3325_n505# a_n3383_n450# 0.101608f
C38 a_1577_n505# a_1777_n450# 0.101608f
C39 a_803_n505# a_745_n450# 0.101608f
C40 a_1261_n450# a_1319_n505# 0.101608f
C41 a_n1319_n450# a_n1061_n450# 0.246592f
C42 a_3125_n505# a_3067_n450# 0.101608f
C43 a_n1061_n450# a_n1261_n505# 0.101608f
C44 a_n2867_n450# a_n3067_n505# 0.101608f
C45 a_n2867_n450# a_n2609_n450# 0.246592f
C46 a_745_n450# a_487_n450# 0.246592f
C47 a_1003_n450# a_1061_n505# 0.101608f
C48 a_n3125_n450# a_n3067_n505# 0.101608f
C49 a_n745_n505# a_n545_n450# 0.101608f
C50 a_n2351_n450# a_n2551_n505# 0.101608f
C51 a_n2035_n505# a_n1835_n450# 0.101608f
C52 a_n287_n450# a_n29_n450# 0.246592f
C53 a_n803_n450# a_n1003_n505# 0.101608f
C54 a_n803_n450# a_n545_n450# 0.246592f
C55 a_n2351_n450# a_n2609_n450# 0.246592f
C56 a_n2093_n450# a_n2293_n505# 0.101608f
C57 a_n2867_n450# a_n2809_n505# 0.101608f
C58 a_1261_n450# a_1003_n450# 0.246592f
C59 a_n1577_n450# a_n1835_n450# 0.246592f
C60 a_2035_n450# a_1835_n505# 0.101608f
C61 a_2035_n450# a_2293_n450# 0.246592f
C62 a_1777_n450# a_1519_n450# 0.246592f
C63 a_229_n450# a_487_n450# 0.246592f
C64 a_2093_n505# a_2293_n450# 0.101608f
C65 a_1519_n450# a_1319_n505# 0.101608f
C66 a_1261_n450# a_1061_n505# 0.101608f
C67 a_1835_n505# a_1777_n450# 0.101608f
C68 a_1003_n450# a_745_n450# 0.246592f
C69 a_2035_n450# a_2093_n505# 0.101608f
C70 a_n287_n450# a_n545_n450# 0.246592f
C71 a_n2093_n450# a_n2351_n450# 0.246592f
C72 a_545_n505# a_745_n450# 0.101608f
C73 a_2867_n505# a_2809_n450# 0.101608f
C74 a_n487_n505# a_n545_n450# 0.101608f
C75 a_n2093_n450# a_n1835_n450# 0.246592f
C76 a_n2609_n450# a_n2551_n505# 0.101608f
C77 a_2035_n450# a_1777_n450# 0.246592f
C78 a_3325_n450# a_n3517_n672# 0.501439f
C79 a_3067_n450# a_n3517_n672# 0.15264f
C80 a_2809_n450# a_n3517_n672# 0.15264f
C81 a_2551_n450# a_n3517_n672# 0.15264f
C82 a_2293_n450# a_n3517_n672# 0.15264f
C83 a_2035_n450# a_n3517_n672# 0.15264f
C84 a_1777_n450# a_n3517_n672# 0.15264f
C85 a_1519_n450# a_n3517_n672# 0.15264f
C86 a_1261_n450# a_n3517_n672# 0.15264f
C87 a_1003_n450# a_n3517_n672# 0.15264f
C88 a_745_n450# a_n3517_n672# 0.15264f
C89 a_487_n450# a_n3517_n672# 0.15264f
C90 a_229_n450# a_n3517_n672# 0.15264f
C91 a_n29_n450# a_n3517_n672# 0.15264f
C92 a_n287_n450# a_n3517_n672# 0.15264f
C93 a_n545_n450# a_n3517_n672# 0.15264f
C94 a_n803_n450# a_n3517_n672# 0.15264f
C95 a_n1061_n450# a_n3517_n672# 0.15264f
C96 a_n1319_n450# a_n3517_n672# 0.15264f
C97 a_n1577_n450# a_n3517_n672# 0.15264f
C98 a_n1835_n450# a_n3517_n672# 0.15264f
C99 a_n2093_n450# a_n3517_n672# 0.15264f
C100 a_n2351_n450# a_n3517_n672# 0.15264f
C101 a_n2609_n450# a_n3517_n672# 0.15264f
C102 a_n2867_n450# a_n3517_n672# 0.15264f
C103 a_n3125_n450# a_n3517_n672# 0.15264f
C104 a_n3383_n450# a_n3517_n672# 0.501439f
C105 a_3125_n505# a_n3517_n672# 0.56045f
C106 a_2867_n505# a_n3517_n672# 0.506278f
C107 a_2609_n505# a_n3517_n672# 0.506278f
C108 a_2351_n505# a_n3517_n672# 0.506278f
C109 a_2093_n505# a_n3517_n672# 0.506278f
C110 a_1835_n505# a_n3517_n672# 0.506278f
C111 a_1577_n505# a_n3517_n672# 0.506278f
C112 a_1319_n505# a_n3517_n672# 0.506278f
C113 a_1061_n505# a_n3517_n672# 0.506278f
C114 a_803_n505# a_n3517_n672# 0.506278f
C115 a_545_n505# a_n3517_n672# 0.506278f
C116 a_287_n505# a_n3517_n672# 0.506278f
C117 a_29_n505# a_n3517_n672# 0.506278f
C118 a_n229_n505# a_n3517_n672# 0.506278f
C119 a_n487_n505# a_n3517_n672# 0.506278f
C120 a_n745_n505# a_n3517_n672# 0.506278f
C121 a_n1003_n505# a_n3517_n672# 0.506278f
C122 a_n1261_n505# a_n3517_n672# 0.506278f
C123 a_n1519_n505# a_n3517_n672# 0.506278f
C124 a_n1777_n505# a_n3517_n672# 0.506278f
C125 a_n2035_n505# a_n3517_n672# 0.506278f
C126 a_n2293_n505# a_n3517_n672# 0.506278f
C127 a_n2551_n505# a_n3517_n672# 0.506278f
C128 a_n2809_n505# a_n3517_n672# 0.506278f
C129 a_n3067_n505# a_n3517_n672# 0.506278f
C130 a_n3325_n505# a_n3517_n672# 0.56045f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_USXRNR a_1448_n255# a_1190_n255# a_358_n200#
+ a_n1648_n255# a_n1706_n200# a_100_n200# a_n674_n200# a_n616_n255# a_n1390_n255#
+ a_674_n255# a_1132_n200# a_n158_n200# a_158_n255# a_616_n200# a_n874_n255# a_n932_n200#
+ a_1648_n200# a_932_n255# a_1390_n200# a_n1448_n200# a_n358_n255# a_n416_n200# a_n1190_n200#
+ a_n1132_n255# a_874_n200# a_416_n255# a_n100_n255# a_n1840_n422#
X0 a_1648_n200# a_1448_n255# a_1390_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X1 a_1132_n200# a_932_n255# a_874_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_874_n200# a_674_n255# a_616_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1390_n200# a_1190_n255# a_1132_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_100_n200# a_n100_n255# a_n158_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n416_n200# a_n616_n255# a_n674_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n158_n200# a_n358_n255# a_n416_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n1448_n200# a_n1648_n255# a_n1706_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X8 a_n1190_n200# a_n1390_n255# a_n1448_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n674_n200# a_n874_n255# a_n932_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n932_n200# a_n1132_n255# a_n1190_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_358_n200# a_158_n255# a_100_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_616_n200# a_416_n255# a_358_n200# a_n1840_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
C0 a_1132_n200# a_1390_n200# 0.110175f
C1 a_n674_n200# a_n416_n200# 0.110175f
C2 a_616_n200# a_874_n200# 0.110175f
C3 a_100_n200# a_n158_n200# 0.110175f
C4 a_n1190_n200# a_n1448_n200# 0.110175f
C5 a_1390_n200# a_1648_n200# 0.110175f
C6 a_n416_n200# a_n158_n200# 0.110175f
C7 a_616_n200# a_358_n200# 0.110175f
C8 a_100_n200# a_358_n200# 0.110175f
C9 a_n1448_n200# a_n1706_n200# 0.110175f
C10 a_n674_n200# a_n932_n200# 0.110175f
C11 a_1132_n200# a_874_n200# 0.110175f
C12 a_n1190_n200# a_n932_n200# 0.110175f
C13 a_1648_n200# a_n1840_n422# 0.241444f
C14 a_n1706_n200# a_n1840_n422# 0.241444f
C15 a_1448_n255# a_n1840_n422# 0.55256f
C16 a_1190_n255# a_n1840_n422# 0.498389f
C17 a_932_n255# a_n1840_n422# 0.498389f
C18 a_674_n255# a_n1840_n422# 0.498389f
C19 a_416_n255# a_n1840_n422# 0.498389f
C20 a_158_n255# a_n1840_n422# 0.498389f
C21 a_n100_n255# a_n1840_n422# 0.498389f
C22 a_n358_n255# a_n1840_n422# 0.498389f
C23 a_n616_n255# a_n1840_n422# 0.498389f
C24 a_n874_n255# a_n1840_n422# 0.498389f
C25 a_n1132_n255# a_n1840_n422# 0.498389f
C26 a_n1390_n255# a_n1840_n422# 0.498389f
C27 a_n1648_n255# a_n1840_n422# 0.55256f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AUMBFF a_n2035_n2564# a_n1519_n2564# a_2035_n2500#
+ a_n1319_n2500# a_1519_n2500# a_n3899_n2500# a_487_n2500# a_545_n2564# a_29_n2564#
+ a_n487_n2564# a_n287_n2500# a_3383_n2564# a_2867_n2564# a_2093_n2564# a_n4099_n2564#
+ a_745_n2500# a_1577_n2564# a_803_n2564# a_n1003_n2564# w_n4615_n2797# a_4099_n2500#
+ a_n545_n2500# a_4157_n2564# a_n745_n2564# a_n3583_n2564# a_1003_n2500# a_n3383_n2500#
+ a_3583_n2500# a_n2867_n2500# a_3641_n2564# a_n2293_n2564# a_2293_n2500# a_n2093_n2500#
+ a_n1777_n2564# a_1777_n2500# a_n29_n2500# a_n1577_n2500# a_n4157_n2500# a_2351_n2564#
+ a_n4357_n2564# a_4357_n2500# a_1835_n2564# a_229_n2500# a_n803_n2500# a_n229_n2564#
+ a_n3841_n2564# a_3841_n2500# a_n3641_n2500# a_1061_n2564# a_n3067_n2564# a_3067_n2500#
+ a_3125_n2564# a_n2551_n2564# a_n2351_n2500# a_2609_n2564# a_2551_n2500# a_n1835_n2500#
+ a_n4415_n2500# a_1319_n2564# a_n1261_n2564# a_1261_n2500# a_n1061_n2500# a_3899_n2564#
+ a_n3125_n2500# a_287_n2564# a_n2809_n2564# a_n3325_n2564# a_3325_n2500# a_n2609_n2500#
+ a_2809_n2500#
X0 a_3067_n2500# a_2867_n2564# a_2809_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X1 a_2809_n2500# a_2609_n2564# a_2551_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X2 a_1777_n2500# a_1577_n2564# a_1519_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X3 a_n4157_n2500# a_n4357_n2564# a_n4415_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=7.25 ps=50.58 w=25 l=1
X4 a_1519_n2500# a_1319_n2564# a_1261_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X5 a_3583_n2500# a_3383_n2564# a_3325_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X6 a_n2867_n2500# a_n3067_n2564# a_n3125_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X7 a_487_n2500# a_287_n2564# a_229_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X8 a_2293_n2500# a_2093_n2564# a_2035_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X9 a_3325_n2500# a_3125_n2564# a_3067_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X10 a_n287_n2500# a_n487_n2564# a_n545_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X11 a_n2609_n2500# a_n2809_n2564# a_n2867_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X12 a_n1577_n2500# a_n1777_n2564# a_n1835_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X13 a_n29_n2500# a_n229_n2564# a_n287_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X14 a_2035_n2500# a_1835_n2564# a_1777_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X15 a_n1319_n2500# a_n1519_n2564# a_n1577_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X16 a_n3383_n2500# a_n3583_n2564# a_n3641_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X17 a_3841_n2500# a_3641_n2564# a_3583_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X18 a_n3125_n2500# a_n3325_n2564# a_n3383_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X19 a_n2093_n2500# a_n2293_n2564# a_n2351_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X20 a_745_n2500# a_545_n2564# a_487_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X21 a_n1835_n2500# a_n2035_n2564# a_n2093_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X22 a_2551_n2500# a_2351_n2564# a_2293_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X23 a_1261_n2500# a_1061_n2564# a_1003_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X24 a_n545_n2500# a_n745_n2564# a_n803_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X25 a_229_n2500# a_29_n2564# a_n29_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X26 a_4099_n2500# a_3899_n2564# a_3841_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X27 a_n3641_n2500# a_n3841_n2564# a_n3899_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X28 a_n2351_n2500# a_n2551_n2564# a_n2609_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X29 a_1003_n2500# a_803_n2564# a_745_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X30 a_n3899_n2500# a_n4099_n2564# a_n4157_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X31 a_n1061_n2500# a_n1261_n2564# a_n1319_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X32 a_n803_n2500# a_n1003_n2564# a_n1061_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=3.625 pd=25.29 as=3.625 ps=25.29 w=25 l=1
X33 a_4357_n2500# a_4157_n2564# a_4099_n2500# w_n4615_n2797# sky130_fd_pr__pfet_g5v0d10v5 ad=7.25 pd=50.58 as=3.625 ps=25.29 w=25 l=1
C0 w_n4615_n2797# a_n3067_n2564# 0.307639f
C1 a_29_n2564# a_n29_n2500# 0.539712f
C2 a_n1061_n2500# a_n803_n2500# 1.36521f
C3 w_n4615_n2797# a_n4099_n2564# 0.307639f
C4 a_3125_n2564# w_n4615_n2797# 0.307639f
C5 a_29_n2564# w_n4615_n2797# 0.307639f
C6 a_n1061_n2500# a_n1003_n2564# 0.539712f
C7 a_n545_n2500# a_n803_n2500# 1.36521f
C8 a_2551_n2500# a_2809_n2500# 1.36521f
C9 w_n4615_n2797# a_3641_n2564# 0.307639f
C10 w_n4615_n2797# a_n4357_n2564# 0.34286f
C11 a_803_n2564# a_745_n2500# 0.539712f
C12 a_545_n2564# a_487_n2500# 0.539712f
C13 a_n1519_n2564# w_n4615_n2797# 0.307639f
C14 a_3383_n2564# a_3325_n2500# 0.539712f
C15 a_n2093_n2500# a_n1835_n2500# 1.36521f
C16 w_n4615_n2797# a_4357_n2500# 1.42757f
C17 a_n1777_n2564# a_n1835_n2500# 0.539712f
C18 a_n2551_n2564# a_n2351_n2500# 0.539712f
C19 a_n4357_n2564# a_n4415_n2500# 0.539712f
C20 w_n4615_n2797# a_1577_n2564# 0.307639f
C21 a_2609_n2564# a_2809_n2500# 0.539712f
C22 a_n287_n2500# a_n29_n2500# 1.36521f
C23 a_n4157_n2500# a_n4415_n2500# 1.36521f
C24 a_2551_n2500# a_2351_n2564# 0.539712f
C25 a_2035_n2500# a_1835_n2564# 0.539712f
C26 a_229_n2500# a_n29_n2500# 1.36521f
C27 a_3067_n2500# a_3125_n2564# 0.539712f
C28 a_1519_n2500# a_1261_n2500# 1.36521f
C29 a_n3583_n2564# a_n3383_n2500# 0.539712f
C30 a_n229_n2564# a_n29_n2500# 0.539712f
C31 a_2351_n2564# a_2293_n2500# 0.539712f
C32 a_n2551_n2564# w_n4615_n2797# 0.307639f
C33 a_4099_n2500# a_4357_n2500# 1.36521f
C34 a_n2809_n2564# a_n2867_n2500# 0.539712f
C35 w_n4615_n2797# a_n229_n2564# 0.307639f
C36 a_2867_n2564# w_n4615_n2797# 0.307639f
C37 w_n4615_n2797# a_2351_n2564# 0.307639f
C38 a_n1261_n2564# w_n4615_n2797# 0.307639f
C39 a_1777_n2500# a_1577_n2564# 0.539712f
C40 a_745_n2500# a_487_n2500# 1.36521f
C41 a_2093_n2564# a_2035_n2500# 0.539712f
C42 a_4099_n2500# a_3841_n2500# 1.36521f
C43 a_n4157_n2500# a_n4099_n2564# 0.539712f
C44 w_n4615_n2797# a_1835_n2564# 0.307639f
C45 w_n4615_n2797# a_287_n2564# 0.307639f
C46 w_n4615_n2797# a_n3325_n2564# 0.307639f
C47 a_3583_n2500# a_3641_n2564# 0.539712f
C48 a_n3125_n2500# a_n3067_n2564# 0.539712f
C49 a_3067_n2500# a_2809_n2500# 1.36521f
C50 a_3899_n2564# w_n4615_n2797# 0.307639f
C51 a_n4157_n2500# a_n4357_n2564# 0.539712f
C52 a_n3125_n2500# a_n3383_n2500# 1.36521f
C53 a_n287_n2500# a_n545_n2500# 1.36521f
C54 a_1319_n2564# a_1519_n2500# 0.539712f
C55 w_n4615_n2797# a_n2035_n2564# 0.307639f
C56 a_2093_n2564# a_2293_n2500# 0.539712f
C57 w_n4615_n2797# a_4157_n2564# 0.34286f
C58 w_n4615_n2797# a_n487_n2564# 0.307639f
C59 a_3067_n2500# a_3325_n2500# 1.36521f
C60 a_1519_n2500# a_1777_n2500# 1.36521f
C61 a_n1061_n2500# a_n1319_n2500# 1.36521f
C62 a_2093_n2564# w_n4615_n2797# 0.307639f
C63 a_n1061_n2500# a_n1261_n2564# 0.539712f
C64 a_n1777_n2564# a_n1577_n2500# 0.539712f
C65 a_1777_n2500# a_1835_n2564# 0.539712f
C66 a_4099_n2500# a_3899_n2564# 0.539712f
C67 a_3125_n2564# a_3325_n2500# 0.539712f
C68 a_n2551_n2564# a_n2609_n2500# 0.539712f
C69 a_1261_n2500# a_1003_n2500# 1.36521f
C70 a_3067_n2500# a_2867_n2564# 0.539712f
C71 a_n2093_n2500# a_n2035_n2564# 0.539712f
C72 a_3583_n2500# a_3841_n2500# 1.36521f
C73 a_n3841_n2564# a_n3899_n2500# 0.539712f
C74 a_n3583_n2564# a_n3641_n2500# 0.539712f
C75 a_2035_n2500# a_2293_n2500# 1.36521f
C76 a_3641_n2564# a_3841_n2500# 0.539712f
C77 a_3325_n2500# a_3583_n2500# 1.36521f
C78 w_n4615_n2797# a_n745_n2564# 0.307639f
C79 a_1061_n2564# a_1003_n2500# 0.539712f
C80 a_29_n2564# a_229_n2500# 0.539712f
C81 a_n3841_n2564# a_n3641_n2500# 0.539712f
C82 a_n2609_n2500# a_n2867_n2500# 1.36521f
C83 a_n2351_n2500# a_n2293_n2564# 0.539712f
C84 a_1061_n2564# a_1261_n2500# 0.539712f
C85 a_4099_n2500# a_4157_n2564# 0.539712f
C86 a_2551_n2500# a_2293_n2500# 1.36521f
C87 a_n3899_n2500# a_n4099_n2564# 0.539712f
C88 a_n3067_n2564# a_n2867_n2500# 0.539712f
C89 a_3383_n2564# w_n4615_n2797# 0.307639f
C90 a_n3641_n2500# a_n3383_n2500# 1.36521f
C91 a_n4157_n2500# a_n3899_n2500# 1.36521f
C92 a_n545_n2500# a_n487_n2564# 0.539712f
C93 a_n745_n2564# a_n803_n2500# 0.539712f
C94 a_2551_n2500# a_2609_n2564# 0.539712f
C95 a_1061_n2564# w_n4615_n2797# 0.307639f
C96 a_229_n2500# a_487_n2500# 1.36521f
C97 a_n3325_n2564# a_n3383_n2500# 0.539712f
C98 w_n4615_n2797# a_n2293_n2564# 0.307639f
C99 w_n4615_n2797# a_n2809_n2564# 0.307639f
C100 a_n2093_n2500# a_n2351_n2500# 1.36521f
C101 a_n1319_n2500# a_n1519_n2564# 0.539712f
C102 a_n1577_n2500# a_n1835_n2500# 1.36521f
C103 a_n3125_n2500# a_n2867_n2500# 1.36521f
C104 a_2035_n2500# a_1777_n2500# 1.36521f
C105 w_n4615_n2797# a_545_n2564# 0.307639f
C106 a_2867_n2564# a_2809_n2500# 0.539712f
C107 a_1319_n2564# a_1261_n2500# 0.539712f
C108 a_n3125_n2500# a_n3325_n2564# 0.539712f
C109 a_n745_n2564# a_n545_n2500# 0.539712f
C110 a_n1835_n2500# a_n2035_n2564# 0.539712f
C111 w_n4615_n2797# a_2609_n2564# 0.307639f
C112 a_287_n2564# a_487_n2500# 0.539712f
C113 a_n2093_n2500# a_n2293_n2564# 0.539712f
C114 a_1519_n2500# a_1577_n2564# 0.539712f
C115 a_n229_n2564# a_n287_n2500# 0.539712f
C116 a_n1519_n2564# a_n1577_n2500# 0.539712f
C117 a_745_n2500# a_1003_n2500# 1.36521f
C118 a_803_n2564# a_1003_n2500# 0.539712f
C119 a_1319_n2564# w_n4615_n2797# 0.307639f
C120 w_n4615_n2797# a_n1777_n2564# 0.307639f
C121 w_n4615_n2797# a_n4415_n2500# 1.42757f
C122 a_n2351_n2500# a_n2609_n2500# 1.36521f
C123 w_n4615_n2797# a_n1003_n2564# 0.307639f
C124 a_3899_n2564# a_3841_n2500# 0.539712f
C125 a_4357_n2500# a_4157_n2564# 0.539712f
C126 a_n1319_n2500# a_n1261_n2564# 0.539712f
C127 a_229_n2500# a_287_n2564# 0.539712f
C128 a_n3641_n2500# a_n3899_n2500# 1.36521f
C129 a_545_n2564# a_745_n2500# 0.539712f
C130 a_803_n2564# w_n4615_n2797# 0.307639f
C131 a_n3583_n2564# w_n4615_n2797# 0.307639f
C132 a_n2809_n2564# a_n2609_n2500# 0.539712f
C133 a_n287_n2500# a_n487_n2564# 0.539712f
C134 a_3383_n2564# a_3583_n2500# 0.539712f
C135 w_n4615_n2797# a_n3841_n2564# 0.307639f
C136 a_n1003_n2564# a_n803_n2500# 0.539712f
C137 a_n1319_n2500# a_n1577_n2500# 1.36521f
C138 a_4357_n2500# 0 1.21504f
C139 a_4099_n2500# 0 0.690385f
C140 a_3841_n2500# 0 0.690385f
C141 a_3583_n2500# 0 0.690385f
C142 a_3325_n2500# 0 0.690385f
C143 a_3067_n2500# 0 0.690385f
C144 a_2809_n2500# 0 0.690385f
C145 a_2551_n2500# 0 0.690385f
C146 a_2293_n2500# 0 0.690385f
C147 a_2035_n2500# 0 0.690385f
C148 a_1777_n2500# 0 0.690385f
C149 a_1519_n2500# 0 0.690385f
C150 a_1261_n2500# 0 0.690385f
C151 a_1003_n2500# 0 0.690385f
C152 a_745_n2500# 0 0.690385f
C153 a_487_n2500# 0 0.690385f
C154 a_229_n2500# 0 0.690385f
C155 a_n29_n2500# 0 0.690385f
C156 a_n287_n2500# 0 0.690385f
C157 a_n545_n2500# 0 0.690385f
C158 a_n803_n2500# 0 0.690385f
C159 a_n1061_n2500# 0 0.690385f
C160 a_n1319_n2500# 0 0.690385f
C161 a_n1577_n2500# 0 0.690385f
C162 a_n1835_n2500# 0 0.690385f
C163 a_n2093_n2500# 0 0.690385f
C164 a_n2351_n2500# 0 0.690385f
C165 a_n2609_n2500# 0 0.690385f
C166 a_n2867_n2500# 0 0.690385f
C167 a_n3125_n2500# 0 0.690385f
C168 a_n3383_n2500# 0 0.690385f
C169 a_n3641_n2500# 0 0.690385f
C170 a_n3899_n2500# 0 0.690385f
C171 a_n4157_n2500# 0 0.690385f
C172 a_n4415_n2500# 0 1.21504f
C173 a_4157_n2564# 0 0.253452f
C174 a_3899_n2564# 0 0.231023f
C175 a_3641_n2564# 0 0.231023f
C176 a_3383_n2564# 0 0.231023f
C177 a_3125_n2564# 0 0.231023f
C178 a_2867_n2564# 0 0.231023f
C179 a_2609_n2564# 0 0.231023f
C180 a_2351_n2564# 0 0.231023f
C181 a_2093_n2564# 0 0.231023f
C182 a_1835_n2564# 0 0.231023f
C183 a_1577_n2564# 0 0.231023f
C184 a_1319_n2564# 0 0.231023f
C185 a_1061_n2564# 0 0.231023f
C186 a_803_n2564# 0 0.231023f
C187 a_545_n2564# 0 0.231023f
C188 a_287_n2564# 0 0.231023f
C189 a_29_n2564# 0 0.231023f
C190 a_n229_n2564# 0 0.231023f
C191 a_n487_n2564# 0 0.231023f
C192 a_n745_n2564# 0 0.231023f
C193 a_n1003_n2564# 0 0.231023f
C194 a_n1261_n2564# 0 0.231023f
C195 a_n1519_n2564# 0 0.231023f
C196 a_n1777_n2564# 0 0.231023f
C197 a_n2035_n2564# 0 0.231023f
C198 a_n2293_n2564# 0 0.231023f
C199 a_n2551_n2564# 0 0.231023f
C200 a_n2809_n2564# 0 0.231023f
C201 a_n3067_n2564# 0 0.231023f
C202 a_n3325_n2564# 0 0.231023f
C203 a_n3583_n2564# 0 0.231023f
C204 a_n3841_n2564# 0 0.231023f
C205 a_n4099_n2564# 0 0.231023f
C206 a_n4357_n2564# 0 0.253452f
C207 w_n4615_n2797# 0 0.163215p
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QL2RRT a_29_n664# a_n1777_n664# a_n2351_n600#
+ a_n745_n664# a_229_n600# a_n1577_n600# a_2867_n664# a_2035_n600# a_803_n664# a_n2035_n664#
+ a_n545_n600# a_3125_n664# a_1835_n664# a_1003_n600# a_n229_n664# w_n3583_n897# a_287_n664#
+ a_n1003_n664# a_n2867_n600# a_3325_n600# a_2093_n664# a_n3325_n664# a_n29_n600#
+ a_487_n600# a_1319_n664# a_2293_n600# a_n3125_n600# a_n2293_n664# a_n1835_n600#
+ a_1061_n664# a_n803_n600# a_1519_n600# a_n2093_n600# a_n1519_n664# a_1261_n600#
+ a_n487_n664# a_n1261_n664# a_2609_n664# a_545_n664# a_n1319_n600# a_n287_n600# a_n1061_n600#
+ a_2351_n664# a_2809_n600# a_1577_n664# a_745_n600# a_n3383_n600# a_n2809_n664# a_2551_n600#
+ a_n2551_n664# a_3067_n600# a_1777_n600# a_n2609_n600# a_n3067_n664#
X0 a_n1835_n600# a_n2035_n664# a_n2093_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_2809_n600# a_2609_n664# a_2551_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2351_n600# a_n2551_n664# a_n2609_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_n2093_n600# a_n2293_n664# a_n2351_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_229_n600# a_29_n664# a_n29_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_n29_n600# a_n229_n664# a_n287_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_3067_n600# a_2867_n664# a_2809_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_n1319_n600# a_n1519_n664# a_n1577_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n545_n600# a_n745_n664# a_n803_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X9 a_2551_n600# a_2351_n664# a_2293_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n3125_n600# a_n3325_n664# a_n3383_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X11 a_n287_n600# a_n487_n664# a_n545_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_2293_n600# a_2093_n664# a_2035_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n2867_n600# a_n3067_n664# a_n3125_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n803_n600# a_n1003_n664# a_n1061_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_n1577_n600# a_n1777_n664# a_n1835_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_1519_n600# a_1319_n664# a_1261_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_n1061_n600# a_n1261_n664# a_n1319_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X18 a_3325_n600# a_3125_n664# a_3067_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X19 a_1003_n600# a_803_n664# a_745_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_487_n600# a_287_n664# a_229_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_745_n600# a_545_n664# a_487_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_2035_n600# a_1835_n664# a_1777_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_n2609_n600# a_n2809_n664# a_n2867_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1777_n600# a_1577_n664# a_1519_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_1261_n600# a_1061_n664# a_1003_n600# w_n3583_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
C0 a_n2609_n600# a_n2809_n664# 0.133664f
C1 a_3125_n664# a_3325_n600# 0.133664f
C2 w_n3583_n897# a_2609_n664# 0.307639f
C3 a_1261_n600# a_1519_n600# 0.328443f
C4 a_1261_n600# a_1003_n600# 0.328443f
C5 a_2609_n664# a_2551_n600# 0.133664f
C6 a_803_n664# a_1003_n600# 0.133664f
C7 a_n1003_n664# a_n803_n600# 0.133664f
C8 w_n3583_n897# a_n1519_n664# 0.307639f
C9 a_1061_n664# a_1003_n600# 0.133664f
C10 w_n3583_n897# a_287_n664# 0.307639f
C11 w_n3583_n897# a_n2551_n664# 0.307639f
C12 a_2093_n664# a_2293_n600# 0.133664f
C13 a_n29_n600# a_n229_n664# 0.133664f
C14 a_n2609_n600# a_n2351_n600# 0.328443f
C15 a_n545_n600# a_n287_n600# 0.328443f
C16 a_803_n664# a_745_n600# 0.133664f
C17 a_n2609_n600# a_n2867_n600# 0.328443f
C18 a_n3383_n600# a_n3325_n664# 0.133664f
C19 a_n1319_n600# a_n1261_n664# 0.133664f
C20 a_n2293_n664# a_n2093_n600# 0.133664f
C21 a_2035_n600# a_1777_n600# 0.328443f
C22 w_n3583_n897# a_n745_n664# 0.307639f
C23 w_n3583_n897# a_29_n664# 0.307639f
C24 a_545_n664# a_487_n600# 0.133664f
C25 a_n545_n600# a_n745_n664# 0.133664f
C26 w_n3583_n897# a_3125_n664# 0.34286f
C27 a_n29_n600# a_n287_n600# 0.328443f
C28 a_3067_n600# a_3325_n600# 0.328443f
C29 a_3067_n600# a_2809_n600# 0.328443f
C30 a_n2035_n664# a_n2093_n600# 0.133664f
C31 w_n3583_n897# a_1319_n664# 0.307639f
C32 w_n3583_n897# a_n3067_n664# 0.307639f
C33 a_2867_n664# a_2809_n600# 0.133664f
C34 w_n3583_n897# a_n1261_n664# 0.307639f
C35 a_745_n600# a_1003_n600# 0.328443f
C36 a_n1319_n600# a_n1061_n600# 0.328443f
C37 w_n3583_n897# a_545_n664# 0.307639f
C38 a_n287_n600# a_n487_n664# 0.133664f
C39 w_n3583_n897# a_1577_n664# 0.307639f
C40 a_1577_n664# a_1777_n600# 0.133664f
C41 a_n2351_n600# a_n2093_n600# 0.328443f
C42 a_n3067_n664# a_n3125_n600# 0.133664f
C43 a_n29_n600# a_29_n664# 0.133664f
C44 w_n3583_n897# a_n2293_n664# 0.307639f
C45 a_229_n600# a_287_n664# 0.133664f
C46 w_n3583_n897# a_n2809_n664# 0.307639f
C47 w_n3583_n897# a_n487_n664# 0.307639f
C48 a_229_n600# a_487_n600# 0.328443f
C49 w_n3583_n897# a_n3325_n664# 0.34286f
C50 a_n2035_n664# a_n1835_n600# 0.133664f
C51 w_n3583_n897# a_n2035_n664# 0.307639f
C52 a_n2551_n664# a_n2351_n600# 0.133664f
C53 a_n1061_n600# a_n1261_n664# 0.133664f
C54 a_n545_n600# a_n487_n664# 0.133664f
C55 w_n3583_n897# a_2867_n664# 0.307639f
C56 w_n3583_n897# a_803_n664# 0.307639f
C57 a_2035_n600# a_1835_n664# 0.133664f
C58 w_n3583_n897# a_2351_n664# 0.307639f
C59 a_n1577_n600# a_n1777_n664# 0.133664f
C60 w_n3583_n897# a_1835_n664# 0.307639f
C61 a_n3325_n664# a_n3125_n600# 0.133664f
C62 w_n3583_n897# a_1061_n664# 0.307639f
C63 a_1777_n600# a_1835_n664# 0.133664f
C64 a_229_n600# a_29_n664# 0.133664f
C65 a_3067_n600# a_3125_n664# 0.133664f
C66 a_2035_n600# a_2293_n600# 0.328443f
C67 a_n745_n664# a_n803_n600# 0.133664f
C68 a_2351_n664# a_2551_n600# 0.133664f
C69 a_1261_n600# a_1319_n664# 0.133664f
C70 w_n3583_n897# a_n1003_n664# 0.307639f
C71 a_n2609_n600# a_n2551_n664# 0.133664f
C72 a_2293_n600# a_2551_n600# 0.328443f
C73 a_2035_n600# a_2093_n664# 0.133664f
C74 a_n545_n600# a_n803_n600# 0.328443f
C75 a_1777_n600# a_1519_n600# 0.328443f
C76 w_n3583_n897# a_2093_n664# 0.307639f
C77 a_745_n600# a_487_n600# 0.328443f
C78 a_n2867_n600# a_n3067_n664# 0.133664f
C79 a_n2867_n600# a_n3125_n600# 0.328443f
C80 a_n29_n600# a_229_n600# 0.328443f
C81 a_2609_n664# a_2809_n600# 0.133664f
C82 a_1319_n664# a_1519_n600# 0.133664f
C83 a_n1519_n664# a_n1577_n600# 0.133664f
C84 a_n1319_n600# a_n1577_n600# 0.328443f
C85 a_n2293_n664# a_n2351_n600# 0.133664f
C86 a_n287_n600# a_n229_n664# 0.133664f
C87 a_n1777_n664# a_n1835_n600# 0.133664f
C88 a_1577_n664# a_1519_n600# 0.133664f
C89 a_n1061_n600# a_n803_n600# 0.328443f
C90 w_n3583_n897# a_n1777_n664# 0.307639f
C91 a_n1061_n600# a_n1003_n664# 0.133664f
C92 a_3067_n600# a_2867_n664# 0.133664f
C93 a_n3383_n600# w_n3583_n897# 0.361553f
C94 a_n2867_n600# a_n2809_n664# 0.133664f
C95 a_n1577_n600# a_n1835_n600# 0.328443f
C96 a_545_n664# a_745_n600# 0.133664f
C97 a_1261_n600# a_1061_n664# 0.133664f
C98 w_n3583_n897# a_3325_n600# 0.361553f
C99 a_n1319_n600# a_n1519_n664# 0.133664f
C100 w_n3583_n897# a_n229_n664# 0.307639f
C101 a_n1835_n600# a_n2093_n600# 0.328443f
C102 a_2809_n600# a_2551_n600# 0.328443f
C103 a_n3383_n600# a_n3125_n600# 0.328443f
C104 a_2293_n600# a_2351_n664# 0.133664f
C105 a_287_n664# a_487_n600# 0.133664f
C106 a_3325_n600# 0 0.298041f
C107 a_3067_n600# 0 0.171485f
C108 a_2809_n600# 0 0.171485f
C109 a_2551_n600# 0 0.171485f
C110 a_2293_n600# 0 0.171485f
C111 a_2035_n600# 0 0.171485f
C112 a_1777_n600# 0 0.171485f
C113 a_1519_n600# 0 0.171485f
C114 a_1261_n600# 0 0.171485f
C115 a_1003_n600# 0 0.171485f
C116 a_745_n600# 0 0.171485f
C117 a_487_n600# 0 0.171485f
C118 a_229_n600# 0 0.171485f
C119 a_n29_n600# 0 0.171485f
C120 a_n287_n600# 0 0.171485f
C121 a_n545_n600# 0 0.171485f
C122 a_n803_n600# 0 0.171485f
C123 a_n1061_n600# 0 0.171485f
C124 a_n1319_n600# 0 0.171485f
C125 a_n1577_n600# 0 0.171485f
C126 a_n1835_n600# 0 0.171485f
C127 a_n2093_n600# 0 0.171485f
C128 a_n2351_n600# 0 0.171485f
C129 a_n2609_n600# 0 0.171485f
C130 a_n2867_n600# 0 0.171485f
C131 a_n3125_n600# 0 0.171485f
C132 a_n3383_n600# 0 0.298041f
C133 a_3125_n664# 0 0.236922f
C134 a_2867_n664# 0 0.214493f
C135 a_2609_n664# 0 0.214493f
C136 a_2351_n664# 0 0.214493f
C137 a_2093_n664# 0 0.214493f
C138 a_1835_n664# 0 0.214493f
C139 a_1577_n664# 0 0.214493f
C140 a_1319_n664# 0 0.214493f
C141 a_1061_n664# 0 0.214493f
C142 a_803_n664# 0 0.214493f
C143 a_545_n664# 0 0.214493f
C144 a_287_n664# 0 0.214493f
C145 a_29_n664# 0 0.214493f
C146 a_n229_n664# 0 0.214493f
C147 a_n487_n664# 0 0.214493f
C148 a_n745_n664# 0 0.214493f
C149 a_n1003_n664# 0 0.214493f
C150 a_n1261_n664# 0 0.214493f
C151 a_n1519_n664# 0 0.214493f
C152 a_n1777_n664# 0 0.214493f
C153 a_n2035_n664# 0 0.214493f
C154 a_n2293_n664# 0 0.214493f
C155 a_n2551_n664# 0 0.214493f
C156 a_n2809_n664# 0 0.214493f
C157 a_n3067_n664# 0 0.214493f
C158 a_n3325_n664# 0 0.236922f
C159 w_n3583_n897# 0 43.5931f
.ends

.subckt sky130_fd_pr__pfet_01v8_U4BBJH a_15_n200# w_n211_n419# a_n33_n297# 0 a_n73_n200#
X0 a_15_n200# a_n33_n297# a_n73_n200# w_n211_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
C0 w_n211_n419# a_n73_n200# 0.142661f
C1 w_n211_n419# a_n33_n297# 0.240434f
C2 w_n211_n419# a_15_n200# 0.142661f
C3 a_15_n200# a_n73_n200# 0.321048f
C4 a_n33_n297# 0 0.119141f
C5 w_n211_n419# 0 1.5811f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QTY6KC a_287_n464# a_n1003_n464# a_487_n400#
+ a_n29_n400# a_1319_n464# w_n1777_n697# a_1061_n464# a_1519_n400# a_n803_n400# a_n1519_n464#
+ a_1261_n400# a_n487_n464# a_n1261_n464# a_n1319_n400# a_545_n464# a_n287_n400# a_n1061_n400#
+ a_745_n400# a_29_n464# a_n745_n464# a_229_n400# a_n1577_n400# a_803_n464# a_n545_n400#
+ a_1003_n400# a_n229_n464#
X0 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X1 a_n545_n400# a_n745_n464# a_n803_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n287_n400# a_n487_n464# a_n545_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_1519_n400# a_1319_n464# a_1261_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X5 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_1003_n400# a_803_n464# a_745_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_487_n400# a_287_n464# a_229_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_745_n400# a_545_n464# a_487_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_1261_n400# a_1061_n464# a_1003_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n29_n400# a_n229_n464# a_n287_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_229_n400# a_29_n464# a_n29_n400# w_n1777_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
C0 w_n1777_n697# a_29_n464# 0.307639f
C1 w_n1777_n697# a_803_n464# 0.307639f
C2 a_745_n400# a_1003_n400# 0.219309f
C3 a_745_n400# a_487_n400# 0.219309f
C4 w_n1777_n697# a_n1261_n464# 0.307639f
C5 a_n29_n400# a_229_n400# 0.219309f
C6 w_n1777_n697# a_287_n464# 0.307639f
C7 a_1519_n400# a_1261_n400# 0.219309f
C8 a_1261_n400# a_1003_n400# 0.219309f
C9 a_n1061_n400# a_n803_n400# 0.219309f
C10 a_n745_n464# w_n1777_n697# 0.307639f
C11 w_n1777_n697# a_n1577_n400# 0.249341f
C12 w_n1777_n697# a_1519_n400# 0.249341f
C13 w_n1777_n697# a_545_n464# 0.307639f
C14 w_n1777_n697# a_n1519_n464# 0.34286f
C15 a_n1319_n400# a_n1577_n400# 0.219309f
C16 w_n1777_n697# a_n229_n464# 0.307639f
C17 w_n1777_n697# a_1319_n464# 0.34286f
C18 a_n1319_n400# a_n1061_n400# 0.219309f
C19 w_n1777_n697# a_1061_n464# 0.307639f
C20 a_n29_n400# a_n287_n400# 0.219309f
C21 a_229_n400# a_487_n400# 0.219309f
C22 a_n287_n400# a_n545_n400# 0.219309f
C23 w_n1777_n697# a_n487_n464# 0.307639f
C24 w_n1777_n697# a_n1003_n464# 0.307639f
C25 a_n545_n400# a_n803_n400# 0.219309f
C26 a_1519_n400# 0 0.201515f
C27 a_1261_n400# 0 0.116864f
C28 a_1003_n400# 0 0.116864f
C29 a_745_n400# 0 0.116864f
C30 a_487_n400# 0 0.116864f
C31 a_229_n400# 0 0.116864f
C32 a_n29_n400# 0 0.116864f
C33 a_n287_n400# 0 0.116864f
C34 a_n545_n400# 0 0.116864f
C35 a_n803_n400# 0 0.116864f
C36 a_n1061_n400# 0 0.116864f
C37 a_n1319_n400# 0 0.116864f
C38 a_n1577_n400# 0 0.201515f
C39 a_1319_n464# 0 0.233871f
C40 a_1061_n464# 0 0.211442f
C41 a_803_n464# 0 0.211442f
C42 a_545_n464# 0 0.211442f
C43 a_287_n464# 0 0.211442f
C44 a_29_n464# 0 0.211442f
C45 a_n229_n464# 0 0.211442f
C46 a_n487_n464# 0 0.211442f
C47 a_n745_n464# 0 0.211442f
C48 a_n1003_n464# 0 0.211442f
C49 a_n1261_n464# 0 0.211442f
C50 a_n1519_n464# 0 0.233871f
C51 w_n1777_n697# 0 17.4861f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z a_1519_n450# a_n803_n450# a_n2093_n450#
+ a_n2551_n505# a_1261_n450# a_29_n505# a_n1777_n505# a_n3067_n505# a_n1319_n450#
+ a_3641_n505# a_3583_n450# a_n4033_n672# a_n287_n450# a_n1061_n450# a_2867_n505#
+ a_n745_n505# a_2809_n450# a_803_n505# a_n2035_n505# a_745_n450# a_n3383_n450# a_n3841_n505#
+ a_2551_n450# a_3125_n505# a_1835_n505# a_3067_n450# a_1777_n450# a_n2609_n450# a_n229_n505#
+ a_n1003_n505# a_n2351_n450# a_287_n505# a_2093_n505# a_229_n450# a_n1577_n450# a_n3325_n505#
+ a_2035_n450# a_3841_n450# a_1319_n505# a_n545_n450# a_n3899_n450# a_1061_n505# a_n2293_n505#
+ a_1003_n450# a_n3641_n450# a_3383_n505# a_n1519_n505# a_n2867_n450# a_n487_n505#
+ a_3325_n450# a_n1261_n505# a_2609_n505# a_n29_n450# a_545_n505# a_487_n450# a_2351_n505#
+ a_n3583_n505# a_2293_n450# a_n1835_n450# a_n3125_n450# a_1577_n505# a_n2809_n505#
X0 a_n2351_n450# a_n2551_n505# a_n2609_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X1 a_n2093_n450# a_n2293_n505# a_n2351_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X2 a_229_n450# a_29_n505# a_n29_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X3 a_n29_n450# a_n229_n505# a_n287_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X4 a_3067_n450# a_2867_n505# a_2809_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X5 a_n1319_n450# a_n1519_n505# a_n1577_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X6 a_n545_n450# a_n745_n505# a_n803_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X7 a_2551_n450# a_2351_n505# a_2293_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X8 a_n3125_n450# a_n3325_n505# a_n3383_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X9 a_n287_n450# a_n487_n505# a_n545_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X10 a_2293_n450# a_2093_n505# a_2035_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X11 a_n2867_n450# a_n3067_n505# a_n3125_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X12 a_n803_n450# a_n1003_n505# a_n1061_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X13 a_n1577_n450# a_n1777_n505# a_n1835_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X14 a_n3641_n450# a_n3841_n505# a_n3899_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=1
X15 a_n3383_n450# a_n3583_n505# a_n3641_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X16 a_1519_n450# a_1319_n505# a_1261_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X17 a_n1061_n450# a_n1261_n505# a_n1319_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X18 a_3325_n450# a_3125_n505# a_3067_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X19 a_1003_n450# a_803_n505# a_745_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X20 a_745_n450# a_545_n505# a_487_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X21 a_487_n450# a_287_n505# a_229_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X22 a_2035_n450# a_1835_n505# a_1777_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X23 a_n2609_n450# a_n2809_n505# a_n2867_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X24 a_1777_n450# a_1577_n505# a_1519_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X25 a_3841_n450# a_3641_n505# a_3583_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=1
X26 a_3583_n450# a_3383_n505# a_3325_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X27 a_1261_n450# a_1061_n505# a_1003_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X28 a_n1835_n450# a_n2035_n505# a_n2093_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
X29 a_2809_n450# a_2609_n505# a_2551_n450# a_n4033_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=1
C0 a_n545_n450# a_n487_n505# 0.101608f
C1 a_n3641_n450# a_n3899_n450# 0.246592f
C2 a_n2093_n450# a_n2351_n450# 0.246592f
C3 a_n1835_n450# a_n1777_n505# 0.101608f
C4 a_487_n450# a_545_n505# 0.101608f
C5 a_n1061_n450# a_n1319_n450# 0.246592f
C6 a_n1519_n505# a_n1319_n450# 0.101608f
C7 a_2035_n450# a_2093_n505# 0.101608f
C8 a_n29_n450# a_229_n450# 0.246592f
C9 a_n1261_n505# a_n1319_n450# 0.101608f
C10 a_2351_n505# a_2551_n450# 0.101608f
C11 a_3383_n505# a_3583_n450# 0.101608f
C12 a_2293_n450# a_2551_n450# 0.246592f
C13 a_1777_n450# a_1577_n505# 0.101608f
C14 a_n2867_n450# a_n3125_n450# 0.246592f
C15 a_n1519_n505# a_n1577_n450# 0.101608f
C16 a_3841_n450# a_3583_n450# 0.246592f
C17 a_n29_n450# a_n229_n505# 0.101608f
C18 a_2351_n505# a_2293_n450# 0.101608f
C19 a_3067_n450# a_2867_n505# 0.101608f
C20 a_1777_n450# a_1519_n450# 0.246592f
C21 a_745_n450# a_1003_n450# 0.246592f
C22 a_745_n450# a_487_n450# 0.246592f
C23 a_3383_n505# a_3325_n450# 0.101608f
C24 a_n3067_n505# a_n3125_n450# 0.101608f
C25 a_n1577_n450# a_n1319_n450# 0.246592f
C26 a_n3641_n450# a_n3383_n450# 0.246592f
C27 a_3067_n450# a_3325_n450# 0.246592f
C28 a_n287_n450# a_n487_n505# 0.101608f
C29 a_1519_n450# a_1319_n505# 0.101608f
C30 a_n803_n450# a_n1003_n505# 0.101608f
C31 a_2609_n505# a_2551_n450# 0.101608f
C32 a_n2609_n450# a_n2351_n450# 0.246592f
C33 a_803_n505# a_1003_n450# 0.101608f
C34 a_3583_n450# a_3325_n450# 0.246592f
C35 a_3841_n450# a_3641_n505# 0.101608f
C36 a_n545_n450# a_n287_n450# 0.246592f
C37 a_3067_n450# a_3125_n505# 0.101608f
C38 a_3641_n505# a_3583_n450# 0.101608f
C39 a_n3067_n505# a_n2867_n450# 0.101608f
C40 a_n2609_n450# a_n2809_n505# 0.101608f
C41 a_1261_n450# a_1003_n450# 0.246592f
C42 a_n3641_n450# a_n3583_n505# 0.101608f
C43 a_n803_n450# a_n745_n505# 0.101608f
C44 a_2809_n450# a_2551_n450# 0.246592f
C45 a_n2093_n450# a_n2293_n505# 0.101608f
C46 a_3067_n450# a_2809_n450# 0.246592f
C47 a_n3325_n505# a_n3383_n450# 0.101608f
C48 a_n1835_n450# a_n1577_n450# 0.246592f
C49 a_1519_n450# a_1261_n450# 0.246592f
C50 a_2035_n450# a_2293_n450# 0.246592f
C51 a_n803_n450# a_n1061_n450# 0.246592f
C52 a_745_n450# a_545_n505# 0.101608f
C53 a_n1061_n450# a_n1003_n505# 0.101608f
C54 a_3125_n505# a_3325_n450# 0.101608f
C55 a_2809_n450# a_2867_n505# 0.101608f
C56 a_1061_n505# a_1261_n450# 0.101608f
C57 a_n3325_n505# a_n3125_n450# 0.101608f
C58 a_n2551_n505# a_n2351_n450# 0.101608f
C59 a_n803_n450# a_n545_n450# 0.246592f
C60 a_n1835_n450# a_n2093_n450# 0.246592f
C61 a_1777_n450# a_1835_n505# 0.101608f
C62 a_2293_n450# a_2093_n505# 0.101608f
C63 a_n2551_n505# a_n2609_n450# 0.101608f
C64 a_n2293_n505# a_n2351_n450# 0.101608f
C65 a_1777_n450# a_2035_n450# 0.246592f
C66 a_29_n505# a_229_n450# 0.101608f
C67 a_n745_n505# a_n545_n450# 0.101608f
C68 a_n3583_n505# a_n3383_n450# 0.101608f
C69 a_n1835_n450# a_n2035_n505# 0.101608f
C70 a_287_n505# a_487_n450# 0.101608f
C71 a_1519_n450# a_1577_n505# 0.101608f
C72 a_2809_n450# a_2609_n505# 0.101608f
C73 a_n2867_n450# a_n2809_n505# 0.101608f
C74 a_29_n505# a_n29_n450# 0.101608f
C75 a_487_n450# a_229_n450# 0.246592f
C76 a_n3383_n450# a_n3125_n450# 0.246592f
C77 a_n2867_n450# a_n2609_n450# 0.246592f
C78 a_n2093_n450# a_n2035_n505# 0.101608f
C79 a_1835_n505# a_2035_n450# 0.101608f
C80 a_n3641_n450# a_n3841_n505# 0.101608f
C81 a_1061_n505# a_1003_n450# 0.101608f
C82 a_n1777_n505# a_n1577_n450# 0.101608f
C83 a_n1061_n450# a_n1261_n505# 0.101608f
C84 a_n29_n450# a_n287_n450# 0.246592f
C85 a_1319_n505# a_1261_n450# 0.101608f
C86 a_n3841_n505# a_n3899_n450# 0.101608f
C87 a_287_n505# a_229_n450# 0.101608f
C88 a_745_n450# a_803_n505# 0.101608f
C89 a_n287_n450# a_n229_n505# 0.101608f
C90 a_3841_n450# a_n4033_n672# 0.501439f
C91 a_3583_n450# a_n4033_n672# 0.15264f
C92 a_3325_n450# a_n4033_n672# 0.15264f
C93 a_3067_n450# a_n4033_n672# 0.15264f
C94 a_2809_n450# a_n4033_n672# 0.15264f
C95 a_2551_n450# a_n4033_n672# 0.15264f
C96 a_2293_n450# a_n4033_n672# 0.15264f
C97 a_2035_n450# a_n4033_n672# 0.15264f
C98 a_1777_n450# a_n4033_n672# 0.15264f
C99 a_1519_n450# a_n4033_n672# 0.15264f
C100 a_1261_n450# a_n4033_n672# 0.15264f
C101 a_1003_n450# a_n4033_n672# 0.15264f
C102 a_745_n450# a_n4033_n672# 0.15264f
C103 a_487_n450# a_n4033_n672# 0.15264f
C104 a_229_n450# a_n4033_n672# 0.15264f
C105 a_n29_n450# a_n4033_n672# 0.15264f
C106 a_n287_n450# a_n4033_n672# 0.15264f
C107 a_n545_n450# a_n4033_n672# 0.15264f
C108 a_n803_n450# a_n4033_n672# 0.15264f
C109 a_n1061_n450# a_n4033_n672# 0.15264f
C110 a_n1319_n450# a_n4033_n672# 0.15264f
C111 a_n1577_n450# a_n4033_n672# 0.15264f
C112 a_n1835_n450# a_n4033_n672# 0.15264f
C113 a_n2093_n450# a_n4033_n672# 0.15264f
C114 a_n2351_n450# a_n4033_n672# 0.15264f
C115 a_n2609_n450# a_n4033_n672# 0.15264f
C116 a_n2867_n450# a_n4033_n672# 0.15264f
C117 a_n3125_n450# a_n4033_n672# 0.15264f
C118 a_n3383_n450# a_n4033_n672# 0.15264f
C119 a_n3641_n450# a_n4033_n672# 0.15264f
C120 a_n3899_n450# a_n4033_n672# 0.501439f
C121 a_3641_n505# a_n4033_n672# 0.56045f
C122 a_3383_n505# a_n4033_n672# 0.506278f
C123 a_3125_n505# a_n4033_n672# 0.506278f
C124 a_2867_n505# a_n4033_n672# 0.506278f
C125 a_2609_n505# a_n4033_n672# 0.506278f
C126 a_2351_n505# a_n4033_n672# 0.506278f
C127 a_2093_n505# a_n4033_n672# 0.506278f
C128 a_1835_n505# a_n4033_n672# 0.506278f
C129 a_1577_n505# a_n4033_n672# 0.506278f
C130 a_1319_n505# a_n4033_n672# 0.506278f
C131 a_1061_n505# a_n4033_n672# 0.506278f
C132 a_803_n505# a_n4033_n672# 0.506278f
C133 a_545_n505# a_n4033_n672# 0.506278f
C134 a_287_n505# a_n4033_n672# 0.506278f
C135 a_29_n505# a_n4033_n672# 0.506278f
C136 a_n229_n505# a_n4033_n672# 0.506278f
C137 a_n487_n505# a_n4033_n672# 0.506278f
C138 a_n745_n505# a_n4033_n672# 0.506278f
C139 a_n1003_n505# a_n4033_n672# 0.506278f
C140 a_n1261_n505# a_n4033_n672# 0.506278f
C141 a_n1519_n505# a_n4033_n672# 0.506278f
C142 a_n1777_n505# a_n4033_n672# 0.506278f
C143 a_n2035_n505# a_n4033_n672# 0.506278f
C144 a_n2293_n505# a_n4033_n672# 0.506278f
C145 a_n2551_n505# a_n4033_n672# 0.506278f
C146 a_n2809_n505# a_n4033_n672# 0.506278f
C147 a_n3067_n505# a_n4033_n672# 0.506278f
C148 a_n3325_n505# a_n4033_n672# 0.506278f
C149 a_n3583_n505# a_n4033_n672# 0.506278f
C150 a_n3841_n505# a_n4033_n672# 0.56045f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QTY6H6 a_1261_n200# a_n487_n264# a_n1261_n264#
+ a_n1319_n200# a_545_n264# a_n287_n200# a_n1061_n200# a_745_n200# a_29_n264# a_229_n200#
+ a_n745_n264# a_n1577_n200# a_803_n264# a_n545_n200# a_1003_n200# a_n229_n264# a_n1003_n264#
+ a_287_n264# a_487_n200# a_n29_n200# a_1319_n264# a_1061_n264# w_n1777_n497# a_n803_n200#
+ a_1519_n200# a_n1519_n264#
X0 a_745_n200# a_545_n264# a_487_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1003_n200# a_803_n264# a_745_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_487_n200# a_287_n264# a_229_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1261_n200# a_1061_n264# a_1003_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n29_n200# a_n229_n264# a_n287_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_229_n200# a_29_n264# a_n29_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n1319_n200# a_n1519_n264# a_n1577_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X7 a_n545_n200# a_n745_n264# a_n803_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n803_n200# a_n1003_n264# a_n1061_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n287_n200# a_n487_n264# a_n545_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_1519_n200# a_1319_n264# a_1261_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X11 a_n1061_n200# a_n1261_n264# a_n1319_n200# w_n1777_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
C0 w_n1777_n497# a_803_n264# 0.307639f
C1 a_n545_n200# a_n803_n200# 0.110175f
C2 w_n1777_n497# a_545_n264# 0.307639f
C3 w_n1777_n497# a_29_n264# 0.307639f
C4 a_n1061_n200# a_n803_n200# 0.110175f
C5 a_1003_n200# a_1261_n200# 0.110175f
C6 a_n29_n200# a_229_n200# 0.110175f
C7 w_n1777_n497# a_1061_n264# 0.307639f
C8 a_n1577_n200# a_n1319_n200# 0.110175f
C9 a_n1519_n264# w_n1777_n497# 0.34286f
C10 a_n745_n264# w_n1777_n497# 0.307639f
C11 w_n1777_n497# a_n1003_n264# 0.307639f
C12 w_n1777_n497# a_n229_n264# 0.307639f
C13 a_n287_n200# a_n545_n200# 0.110175f
C14 a_n287_n200# a_n29_n200# 0.110175f
C15 a_n1061_n200# a_n1319_n200# 0.110175f
C16 w_n1777_n497# a_1319_n264# 0.34286f
C17 w_n1777_n497# a_n1261_n264# 0.307639f
C18 a_1003_n200# a_745_n200# 0.110175f
C19 a_1261_n200# a_1519_n200# 0.110175f
C20 a_287_n264# w_n1777_n497# 0.307639f
C21 a_745_n200# a_487_n200# 0.110175f
C22 w_n1777_n497# a_n1577_n200# 0.137129f
C23 a_487_n200# a_229_n200# 0.110175f
C24 w_n1777_n497# a_1519_n200# 0.137129f
C25 w_n1777_n497# a_n487_n264# 0.307639f
C26 a_1519_n200# 0 0.104989f
C27 a_n1577_n200# 0 0.104989f
C28 a_1319_n264# 0 0.227252f
C29 a_1061_n264# 0 0.204823f
C30 a_803_n264# 0 0.204823f
C31 a_545_n264# 0 0.204823f
C32 a_287_n264# 0 0.204823f
C33 a_29_n264# 0 0.204823f
C34 a_n229_n264# 0 0.204823f
C35 a_n487_n264# 0 0.204823f
C36 a_n745_n264# 0 0.204823f
C37 a_n1003_n264# 0 0.204823f
C38 a_n1261_n264# 0 0.204823f
C39 a_n1519_n264# 0 0.227252f
C40 w_n1777_n497# 0 12.9886f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_U73S5M a_229_n1000# a_n803_n1000# a_545_n1055#
+ a_29_n1055# a_n487_n1055# a_n4549_n1222# a_n3641_n1000# a_3841_n1000# a_3067_n1000#
+ a_3383_n1055# a_2867_n1055# a_2551_n1000# a_n2351_n1000# a_n1835_n1000# a_n4415_n1000#
+ a_2093_n1055# a_n4099_n1055# a_1577_n1055# a_803_n1055# a_n745_n1055# a_n1003_n1055#
+ a_n1061_n1000# a_4157_n1055# a_n3583_n1055# a_1261_n1000# a_n3125_n1000# a_3641_n1055#
+ a_3325_n1000# a_2809_n1000# a_n2609_n1000# a_n2293_n1055# a_n1777_n1055# a_2035_n1000#
+ a_2351_n1055# a_n4357_n1055# a_1519_n1000# a_n1319_n1000# a_n3899_n1000# a_1835_n1055#
+ a_487_n1000# a_n229_n1055# a_n3841_n1055# a_n287_n1000# a_1061_n1055# a_n3067_n1055#
+ a_3125_n1055# a_n2551_n1055# a_2609_n1055# a_1319_n1055# a_n1261_n1055# a_4099_n1000#
+ a_745_n1000# a_3899_n1055# a_1003_n1000# a_n545_n1000# a_287_n1055# a_n2809_n1055#
+ a_n3325_n1055# a_3583_n1000# a_n3383_n1000# a_n2867_n1000# a_n2035_n1055# a_n2093_n1000#
+ a_n1519_n1055# a_2293_n1000# a_n1577_n1000# a_4357_n1000# a_1777_n1000# a_n29_n1000#
+ a_n4157_n1000#
X0 a_3067_n1000# a_2867_n1055# a_2809_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X1 a_n1319_n1000# a_n1519_n1055# a_n1577_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X2 a_n545_n1000# a_n745_n1055# a_n803_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X3 a_2293_n1000# a_2093_n1055# a_2035_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X4 a_2551_n1000# a_2351_n1055# a_2293_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X5 a_n3125_n1000# a_n3325_n1055# a_n3383_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X6 a_n2867_n1000# a_n3067_n1055# a_n3125_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X7 a_n803_n1000# a_n1003_n1055# a_n1061_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X8 a_n287_n1000# a_n487_n1055# a_n545_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X9 a_n3641_n1000# a_n3841_n1055# a_n3899_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X10 a_n1577_n1000# a_n1777_n1055# a_n1835_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X11 a_1519_n1000# a_1319_n1055# a_1261_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X12 a_n3383_n1000# a_n3583_n1055# a_n3641_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X13 a_3325_n1000# a_3125_n1055# a_3067_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X14 a_n1061_n1000# a_n1261_n1055# a_n1319_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X15 a_745_n1000# a_545_n1055# a_487_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X16 a_1003_n1000# a_803_n1055# a_745_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X17 a_487_n1000# a_287_n1055# a_229_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X18 a_2035_n1000# a_1835_n1055# a_1777_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X19 a_4099_n1000# a_3899_n1055# a_3841_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X20 a_n2609_n1000# a_n2809_n1055# a_n2867_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X21 a_1777_n1000# a_1577_n1055# a_1519_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X22 a_3841_n1000# a_3641_n1055# a_3583_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X23 a_1261_n1000# a_1061_n1055# a_1003_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X24 a_3583_n1000# a_3383_n1055# a_3325_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X25 a_n4157_n1000# a_n4357_n1055# a_n4415_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=2.9 ps=20.58 w=10 l=1
X26 a_n3899_n1000# a_n4099_n1055# a_n4157_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X27 a_n1835_n1000# a_n2035_n1055# a_n2093_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X28 a_2809_n1000# a_2609_n1055# a_2551_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X29 a_n2351_n1000# a_n2551_n1055# a_n2609_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X30 a_4357_n1000# a_4157_n1055# a_4099_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=2.9 pd=20.58 as=1.45 ps=10.29 w=10 l=1
X31 a_n2093_n1000# a_n2293_n1055# a_n2351_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X32 a_n29_n1000# a_n229_n1055# a_n287_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
X33 a_229_n1000# a_29_n1055# a_n29_n1000# a_n4549_n1222# sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.29 as=1.45 ps=10.29 w=10 l=1
C0 a_2351_n1055# a_2551_n1000# 0.219148f
C1 a_n1261_n1055# a_n1319_n1000# 0.219148f
C2 a_487_n1000# a_287_n1055# 0.219148f
C3 a_4099_n1000# a_3899_n1055# 0.219148f
C4 a_n3383_n1000# a_n3583_n1055# 0.219148f
C5 a_n2609_n1000# a_n2867_n1000# 0.54671f
C6 a_n2609_n1000# a_n2551_n1055# 0.219148f
C7 a_n1777_n1055# a_n1835_n1000# 0.219148f
C8 a_3325_n1000# a_3067_n1000# 0.54671f
C9 a_n1577_n1000# a_n1319_n1000# 0.54671f
C10 a_2035_n1000# a_1777_n1000# 0.54671f
C11 a_3583_n1000# a_3641_n1055# 0.219148f
C12 a_n4157_n1000# a_n4357_n1055# 0.219148f
C13 a_n1003_n1055# a_n1061_n1000# 0.219148f
C14 a_n3841_n1055# a_n3641_n1000# 0.219148f
C15 a_1003_n1000# a_745_n1000# 0.54671f
C16 a_3841_n1000# a_3899_n1055# 0.219148f
C17 a_2293_n1000# a_2035_n1000# 0.54671f
C18 a_n29_n1000# a_29_n1055# 0.219148f
C19 a_4357_n1000# a_4157_n1055# 0.219148f
C20 a_1835_n1055# a_1777_n1000# 0.219148f
C21 a_545_n1055# a_745_n1000# 0.219148f
C22 a_3583_n1000# a_3383_n1055# 0.219148f
C23 a_n2035_n1055# a_n1835_n1000# 0.219148f
C24 a_n745_n1055# a_n545_n1000# 0.219148f
C25 a_2809_n1000# a_2609_n1055# 0.219148f
C26 a_229_n1000# a_n29_n1000# 0.54671f
C27 a_3325_n1000# a_3125_n1055# 0.219148f
C28 a_1519_n1000# a_1777_n1000# 0.54671f
C29 a_n803_n1000# a_n545_n1000# 0.54671f
C30 a_n1577_n1000# a_n1777_n1055# 0.219148f
C31 a_n2293_n1055# a_n2351_n1000# 0.219148f
C32 a_1577_n1055# a_1519_n1000# 0.219148f
C33 a_n803_n1000# a_n1061_n1000# 0.54671f
C34 a_1261_n1000# a_1061_n1055# 0.219148f
C35 a_n4157_n1000# a_n4099_n1055# 0.219148f
C36 a_n3125_n1000# a_n2867_n1000# 0.54671f
C37 a_1835_n1055# a_2035_n1000# 0.219148f
C38 a_2867_n1055# a_2809_n1000# 0.219148f
C39 a_n3383_n1000# a_n3641_n1000# 0.54671f
C40 a_n487_n1055# a_n287_n1000# 0.219148f
C41 a_2809_n1000# a_3067_n1000# 0.54671f
C42 a_n1319_n1000# a_n1519_n1055# 0.219148f
C43 a_4099_n1000# a_3841_n1000# 0.54671f
C44 a_3383_n1055# a_3325_n1000# 0.219148f
C45 a_n2093_n1000# a_n1835_n1000# 0.54671f
C46 a_1319_n1055# a_1519_n1000# 0.219148f
C47 a_3583_n1000# a_3325_n1000# 0.54671f
C48 a_1003_n1000# a_803_n1055# 0.219148f
C49 a_n287_n1000# a_n545_n1000# 0.54671f
C50 a_n1577_n1000# a_n1519_n1055# 0.219148f
C51 a_n3067_n1055# a_n2867_n1000# 0.219148f
C52 a_229_n1000# a_29_n1055# 0.219148f
C53 a_n2609_n1000# a_n2809_n1055# 0.219148f
C54 a_1003_n1000# a_1261_n1000# 0.54671f
C55 a_n4415_n1000# a_n4357_n1055# 0.219148f
C56 a_803_n1055# a_745_n1000# 0.219148f
C57 a_n3383_n1000# a_n3125_n1000# 0.54671f
C58 a_2293_n1000# a_2093_n1055# 0.219148f
C59 a_n229_n1055# a_n287_n1000# 0.219148f
C60 a_487_n1000# a_545_n1055# 0.219148f
C61 a_2035_n1000# a_2093_n1055# 0.219148f
C62 a_4099_n1000# a_4157_n1055# 0.219148f
C63 a_2867_n1055# a_3067_n1000# 0.219148f
C64 a_2293_n1000# a_2351_n1055# 0.219148f
C65 a_n29_n1000# a_n287_n1000# 0.54671f
C66 a_1261_n1000# a_1319_n1055# 0.219148f
C67 a_n3067_n1055# a_n3125_n1000# 0.219148f
C68 a_2809_n1000# a_2551_n1000# 0.54671f
C69 a_2293_n1000# a_2551_n1000# 0.54671f
C70 a_n487_n1055# a_n545_n1000# 0.219148f
C71 a_487_n1000# a_745_n1000# 0.54671f
C72 a_n2351_n1000# a_n2609_n1000# 0.54671f
C73 a_n2293_n1055# a_n2093_n1000# 0.219148f
C74 a_n2809_n1055# a_n2867_n1000# 0.219148f
C75 a_n2351_n1000# a_n2093_n1000# 0.54671f
C76 a_2551_n1000# a_2609_n1055# 0.219148f
C77 a_n3899_n1000# a_n4099_n1055# 0.219148f
C78 a_n3641_n1000# a_n3899_n1000# 0.54671f
C79 a_3841_n1000# a_3641_n1055# 0.219148f
C80 a_1261_n1000# a_1519_n1000# 0.54671f
C81 a_n803_n1000# a_n1003_n1055# 0.219148f
C82 a_n3641_n1000# a_n3583_n1055# 0.219148f
C83 a_229_n1000# a_487_n1000# 0.54671f
C84 a_n2351_n1000# a_n2551_n1055# 0.219148f
C85 a_3067_n1000# a_3125_n1055# 0.219148f
C86 a_229_n1000# a_287_n1055# 0.219148f
C87 a_n3841_n1055# a_n3899_n1000# 0.219148f
C88 a_n803_n1000# a_n745_n1055# 0.219148f
C89 a_n1261_n1055# a_n1061_n1000# 0.219148f
C90 a_n1061_n1000# a_n1319_n1000# 0.54671f
C91 a_n3125_n1000# a_n3325_n1055# 0.219148f
C92 a_4099_n1000# a_4357_n1000# 0.54671f
C93 a_1003_n1000# a_1061_n1055# 0.219148f
C94 a_3583_n1000# a_3841_n1000# 0.54671f
C95 a_n2035_n1055# a_n2093_n1000# 0.219148f
C96 a_n4157_n1000# a_n4415_n1000# 0.54671f
C97 a_n229_n1055# a_n29_n1000# 0.219148f
C98 a_n1577_n1000# a_n1835_n1000# 0.54671f
C99 a_n3383_n1000# a_n3325_n1055# 0.219148f
C100 a_1577_n1055# a_1777_n1000# 0.219148f
C101 a_n4157_n1000# a_n3899_n1000# 0.54671f
C102 a_4357_n1000# a_n4549_n1222# 1.07343f
C103 a_4099_n1000# a_n4549_n1222# 0.302848f
C104 a_3841_n1000# a_n4549_n1222# 0.302848f
C105 a_3583_n1000# a_n4549_n1222# 0.302848f
C106 a_3325_n1000# a_n4549_n1222# 0.302848f
C107 a_3067_n1000# a_n4549_n1222# 0.302848f
C108 a_2809_n1000# a_n4549_n1222# 0.302848f
C109 a_2551_n1000# a_n4549_n1222# 0.302848f
C110 a_2293_n1000# a_n4549_n1222# 0.302848f
C111 a_2035_n1000# a_n4549_n1222# 0.302848f
C112 a_1777_n1000# a_n4549_n1222# 0.302848f
C113 a_1519_n1000# a_n4549_n1222# 0.302848f
C114 a_1261_n1000# a_n4549_n1222# 0.302848f
C115 a_1003_n1000# a_n4549_n1222# 0.302848f
C116 a_745_n1000# a_n4549_n1222# 0.302848f
C117 a_487_n1000# a_n4549_n1222# 0.302848f
C118 a_229_n1000# a_n4549_n1222# 0.302848f
C119 a_n29_n1000# a_n4549_n1222# 0.302848f
C120 a_n287_n1000# a_n4549_n1222# 0.302848f
C121 a_n545_n1000# a_n4549_n1222# 0.302848f
C122 a_n803_n1000# a_n4549_n1222# 0.302848f
C123 a_n1061_n1000# a_n4549_n1222# 0.302848f
C124 a_n1319_n1000# a_n4549_n1222# 0.302848f
C125 a_n1577_n1000# a_n4549_n1222# 0.302848f
C126 a_n1835_n1000# a_n4549_n1222# 0.302848f
C127 a_n2093_n1000# a_n4549_n1222# 0.302848f
C128 a_n2351_n1000# a_n4549_n1222# 0.302848f
C129 a_n2609_n1000# a_n4549_n1222# 0.302848f
C130 a_n2867_n1000# a_n4549_n1222# 0.302848f
C131 a_n3125_n1000# a_n4549_n1222# 0.302848f
C132 a_n3383_n1000# a_n4549_n1222# 0.302848f
C133 a_n3641_n1000# a_n4549_n1222# 0.302848f
C134 a_n3899_n1000# a_n4549_n1222# 0.302848f
C135 a_n4157_n1000# a_n4549_n1222# 0.302848f
C136 a_n4415_n1000# a_n4549_n1222# 1.07343f
C137 a_4157_n1055# a_n4549_n1222# 0.579228f
C138 a_3899_n1055# a_n4549_n1222# 0.525056f
C139 a_3641_n1055# a_n4549_n1222# 0.525056f
C140 a_3383_n1055# a_n4549_n1222# 0.525056f
C141 a_3125_n1055# a_n4549_n1222# 0.525056f
C142 a_2867_n1055# a_n4549_n1222# 0.525056f
C143 a_2609_n1055# a_n4549_n1222# 0.525056f
C144 a_2351_n1055# a_n4549_n1222# 0.525056f
C145 a_2093_n1055# a_n4549_n1222# 0.525056f
C146 a_1835_n1055# a_n4549_n1222# 0.525056f
C147 a_1577_n1055# a_n4549_n1222# 0.525056f
C148 a_1319_n1055# a_n4549_n1222# 0.525056f
C149 a_1061_n1055# a_n4549_n1222# 0.525056f
C150 a_803_n1055# a_n4549_n1222# 0.525056f
C151 a_545_n1055# a_n4549_n1222# 0.525056f
C152 a_287_n1055# a_n4549_n1222# 0.525056f
C153 a_29_n1055# a_n4549_n1222# 0.525056f
C154 a_n229_n1055# a_n4549_n1222# 0.525056f
C155 a_n487_n1055# a_n4549_n1222# 0.525056f
C156 a_n745_n1055# a_n4549_n1222# 0.525056f
C157 a_n1003_n1055# a_n4549_n1222# 0.525056f
C158 a_n1261_n1055# a_n4549_n1222# 0.525056f
C159 a_n1519_n1055# a_n4549_n1222# 0.525056f
C160 a_n1777_n1055# a_n4549_n1222# 0.525056f
C161 a_n2035_n1055# a_n4549_n1222# 0.525056f
C162 a_n2293_n1055# a_n4549_n1222# 0.525056f
C163 a_n2551_n1055# a_n4549_n1222# 0.525056f
C164 a_n2809_n1055# a_n4549_n1222# 0.525056f
C165 a_n3067_n1055# a_n4549_n1222# 0.525056f
C166 a_n3325_n1055# a_n4549_n1222# 0.525056f
C167 a_n3583_n1055# a_n4549_n1222# 0.525056f
C168 a_n3841_n1055# a_n4549_n1222# 0.525056f
C169 a_n4099_n1055# a_n4549_n1222# 0.525056f
C170 a_n4357_n1055# a_n4549_n1222# 0.579228f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_PP2RNK a_29_n964# a_n2351_n900# a_229_n900# a_2867_n964#
+ a_n745_n964# a_n1577_n900# a_2035_n900# a_803_n964# a_n2035_n964# a_n545_n900# w_n3325_n1197#
+ a_1835_n964# a_1003_n900# a_n229_n964# a_n1003_n964# a_287_n964# a_n2867_n900# a_2093_n964#
+ a_487_n900# a_n29_n900# a_2293_n900# a_n3125_n900# a_1319_n964# a_n1835_n900# a_1061_n964#
+ a_n2293_n964# a_n803_n900# a_1519_n900# a_n2093_n900# a_n1519_n964# a_1261_n900#
+ a_n487_n964# a_n1261_n964# a_2609_n964# a_n1319_n900# a_545_n964# a_n287_n900# a_2351_n964#
+ a_n1061_n900# a_1577_n964# a_2809_n900# a_745_n900# a_n2809_n964# a_2551_n900# a_n2551_n964#
+ a_3067_n900# a_1777_n900# a_n2609_n900# a_n1777_n964# a_n3067_n964#
X0 a_n2609_n900# a_n2809_n964# a_n2867_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X1 a_1261_n900# a_1061_n964# a_1003_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X2 a_n1835_n900# a_n2035_n964# a_n2093_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X3 a_2809_n900# a_2609_n964# a_2551_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X4 a_n2351_n900# a_n2551_n964# a_n2609_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 a_n2093_n900# a_n2293_n964# a_n2351_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 a_n29_n900# a_n229_n964# a_n287_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X7 a_229_n900# a_29_n964# a_n29_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 a_3067_n900# a_2867_n964# a_2809_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X9 a_n1319_n900# a_n1519_n964# a_n1577_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 a_2551_n900# a_2351_n964# a_2293_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X11 a_n545_n900# a_n745_n964# a_n803_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 a_n287_n900# a_n487_n964# a_n545_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X13 a_2293_n900# a_2093_n964# a_2035_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X14 a_n2867_n900# a_n3067_n964# a_n3125_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X15 a_n803_n900# a_n1003_n964# a_n1061_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X16 a_n1577_n900# a_n1777_n964# a_n1835_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 a_1519_n900# a_1319_n964# a_1261_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X18 a_n1061_n900# a_n1261_n964# a_n1319_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X19 a_1003_n900# a_803_n964# a_745_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X20 a_745_n900# a_545_n964# a_487_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X21 a_487_n900# a_287_n964# a_229_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X22 a_1777_n900# a_1577_n964# a_1519_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X23 a_2035_n900# a_1835_n964# a_1777_n900# w_n3325_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
C0 a_n2035_n964# w_n3325_n1197# 0.307639f
C1 a_n287_n900# a_n29_n900# 0.492143f
C2 a_n487_n964# a_n287_n900# 0.197777f
C3 a_n1319_n900# a_n1261_n964# 0.197777f
C4 a_n287_n900# a_n545_n900# 0.492143f
C5 a_n3125_n900# w_n3325_n1197# 0.529871f
C6 a_n2351_n900# a_n2551_n964# 0.197777f
C7 a_n3067_n964# w_n3325_n1197# 0.34286f
C8 a_2035_n900# a_1777_n900# 0.492143f
C9 a_1835_n964# a_1777_n900# 0.197777f
C10 w_n3325_n1197# a_n1519_n964# 0.307639f
C11 a_2093_n964# w_n3325_n1197# 0.307639f
C12 a_n2609_n900# a_n2809_n964# 0.197777f
C13 a_1319_n964# w_n3325_n1197# 0.307639f
C14 a_n1003_n964# a_n1061_n900# 0.197777f
C15 a_1577_n964# a_1777_n900# 0.197777f
C16 a_1261_n900# a_1519_n900# 0.492143f
C17 a_1319_n964# a_1261_n900# 0.197777f
C18 a_n803_n900# a_n1003_n964# 0.197777f
C19 a_803_n964# a_1003_n900# 0.197777f
C20 a_n1003_n964# w_n3325_n1197# 0.307639f
C21 a_n1577_n900# a_n1519_n964# 0.197777f
C22 a_1835_n964# w_n3325_n1197# 0.307639f
C23 a_n1319_n900# a_n1519_n964# 0.197777f
C24 a_229_n900# a_29_n964# 0.197777f
C25 a_n2351_n900# a_n2609_n900# 0.492143f
C26 a_2293_n900# a_2551_n900# 0.492143f
C27 a_2867_n964# a_2809_n900# 0.197777f
C28 a_n1835_n900# a_n1577_n900# 0.492143f
C29 a_1577_n964# w_n3325_n1197# 0.307639f
C30 a_n1777_n964# w_n3325_n1197# 0.307639f
C31 a_29_n964# w_n3325_n1197# 0.307639f
C32 a_n2293_n964# w_n3325_n1197# 0.307639f
C33 a_229_n900# a_487_n900# 0.492143f
C34 w_n3325_n1197# a_n229_n964# 0.307639f
C35 a_n803_n900# a_n1061_n900# 0.492143f
C36 a_1261_n900# a_1003_n900# 0.492143f
C37 a_n2035_n964# a_n2093_n900# 0.197777f
C38 a_2867_n964# w_n3325_n1197# 0.34286f
C39 a_803_n964# w_n3325_n1197# 0.307639f
C40 a_n2351_n900# a_n2093_n900# 0.492143f
C41 a_2867_n964# a_3067_n900# 0.197777f
C42 a_n1777_n964# a_n1577_n900# 0.197777f
C43 a_n745_n964# a_n803_n900# 0.197777f
C44 a_2809_n900# a_3067_n900# 0.492143f
C45 a_n2551_n964# w_n3325_n1197# 0.307639f
C46 a_2293_n900# a_2351_n964# 0.197777f
C47 a_n3125_n900# a_n3067_n964# 0.197777f
C48 a_2551_n900# a_2809_n900# 0.492143f
C49 a_29_n964# a_n29_n900# 0.197777f
C50 a_n745_n964# w_n3325_n1197# 0.307639f
C51 a_1061_n964# a_1003_n900# 0.197777f
C52 a_n29_n900# a_n229_n964# 0.197777f
C53 a_n1835_n900# a_n2093_n900# 0.492143f
C54 a_1003_n900# a_745_n900# 0.492143f
C55 a_287_n964# a_487_n900# 0.197777f
C56 a_2609_n964# a_2809_n900# 0.197777f
C57 a_545_n964# a_487_n900# 0.197777f
C58 a_287_n964# a_229_n900# 0.197777f
C59 a_3067_n900# w_n3325_n1197# 0.529871f
C60 a_n2035_n964# a_n1835_n900# 0.197777f
C61 a_n1319_n900# a_n1061_n900# 0.492143f
C62 a_229_n900# a_n29_n900# 0.492143f
C63 a_803_n964# a_745_n900# 0.197777f
C64 a_1319_n964# a_1519_n900# 0.197777f
C65 a_287_n964# w_n3325_n1197# 0.307639f
C66 a_n2609_n900# a_n2867_n900# 0.492143f
C67 a_n287_n900# a_n229_n964# 0.197777f
C68 a_745_n900# a_487_n900# 0.492143f
C69 a_n803_n900# a_n545_n900# 0.492143f
C70 a_545_n964# w_n3325_n1197# 0.307639f
C71 a_2609_n964# w_n3325_n1197# 0.307639f
C72 a_n745_n964# a_n545_n900# 0.197777f
C73 a_n487_n964# w_n3325_n1197# 0.307639f
C74 a_n1061_n900# a_n1261_n964# 0.197777f
C75 a_n2609_n900# a_n2551_n964# 0.197777f
C76 a_2293_n900# a_2093_n964# 0.197777f
C77 a_n2293_n964# a_n2093_n900# 0.197777f
C78 a_1061_n964# w_n3325_n1197# 0.307639f
C79 a_n2809_n964# a_n2867_n900# 0.197777f
C80 a_2093_n964# a_2035_n900# 0.197777f
C81 a_2551_n900# a_2609_n964# 0.197777f
C82 a_n1261_n964# w_n3325_n1197# 0.307639f
C83 a_1061_n964# a_1261_n900# 0.197777f
C84 w_n3325_n1197# a_2351_n964# 0.307639f
C85 a_1577_n964# a_1519_n900# 0.197777f
C86 a_n2809_n964# w_n3325_n1197# 0.307639f
C87 a_n2351_n900# a_n2293_n964# 0.197777f
C88 a_n1319_n900# a_n1577_n900# 0.492143f
C89 a_n487_n964# a_n545_n900# 0.197777f
C90 a_2293_n900# a_2035_n900# 0.492143f
C91 a_1777_n900# a_1519_n900# 0.492143f
C92 a_2551_n900# a_2351_n964# 0.197777f
C93 a_n3125_n900# a_n2867_n900# 0.492143f
C94 a_n2867_n900# a_n3067_n964# 0.197777f
C95 a_545_n964# a_745_n900# 0.197777f
C96 a_n1777_n964# a_n1835_n900# 0.197777f
C97 a_2035_n900# a_1835_n964# 0.197777f
C98 a_3067_n900# 0 0.442831f
C99 a_2809_n900# 0 0.253417f
C100 a_2551_n900# 0 0.253417f
C101 a_2293_n900# 0 0.253417f
C102 a_2035_n900# 0 0.253417f
C103 a_1777_n900# 0 0.253417f
C104 a_1519_n900# 0 0.253417f
C105 a_1261_n900# 0 0.253417f
C106 a_1003_n900# 0 0.253417f
C107 a_745_n900# 0 0.253417f
C108 a_487_n900# 0 0.253417f
C109 a_229_n900# 0 0.253417f
C110 a_n29_n900# 0 0.253417f
C111 a_n287_n900# 0 0.253417f
C112 a_n545_n900# 0 0.253417f
C113 a_n803_n900# 0 0.253417f
C114 a_n1061_n900# 0 0.253417f
C115 a_n1319_n900# 0 0.253417f
C116 a_n1577_n900# 0 0.253417f
C117 a_n1835_n900# 0 0.253417f
C118 a_n2093_n900# 0 0.253417f
C119 a_n2351_n900# 0 0.253417f
C120 a_n2609_n900# 0 0.253417f
C121 a_n2867_n900# 0 0.253417f
C122 a_n3125_n900# 0 0.442831f
C123 a_2867_n964# 0 0.253452f
C124 a_2609_n964# 0 0.231023f
C125 a_2351_n964# 0 0.231023f
C126 a_2093_n964# 0 0.231023f
C127 a_1835_n964# 0 0.231023f
C128 a_1577_n964# 0 0.231023f
C129 a_1319_n964# 0 0.231023f
C130 a_1061_n964# 0 0.231023f
C131 a_803_n964# 0 0.231023f
C132 a_545_n964# 0 0.231023f
C133 a_287_n964# 0 0.231023f
C134 a_29_n964# 0 0.231023f
C135 a_n229_n964# 0 0.231023f
C136 a_n487_n964# 0 0.231023f
C137 a_n745_n964# 0 0.231023f
C138 a_n1003_n964# 0 0.231023f
C139 a_n1261_n964# 0 0.231023f
C140 a_n1519_n964# 0 0.231023f
C141 a_n1777_n964# 0 0.231023f
C142 a_n2035_n964# 0 0.231023f
C143 a_n2293_n964# 0 0.231023f
C144 a_n2551_n964# 0 0.231023f
C145 a_n2809_n964# 0 0.231023f
C146 a_n3067_n964# 0 0.253452f
C147 w_n3325_n1197# 0 52.879303f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_79TVLH a_3067_n300# a_1777_n300# a_n2609_n300#
+ a_1061_n355# a_n2293_n355# a_n2351_n300# a_229_n300# a_n1577_n300# a_n1519_n355#
+ a_2035_n300# a_n487_n355# a_n545_n300# a_n1261_n355# a_2609_n355# a_545_n355# a_n3517_n522#
+ a_2351_n355# a_1003_n300# a_1577_n355# a_n2867_n300# a_n2809_n355# a_3325_n300#
+ a_n2551_n355# a_487_n300# a_n29_n300# a_n3067_n355# a_29_n355# a_n1777_n355# a_2293_n300#
+ a_n1835_n300# a_n3125_n300# a_n745_n355# a_2867_n355# a_1519_n300# a_n803_n300#
+ a_n2093_n300# a_803_n355# a_n2035_n355# a_1261_n300# a_n1319_n300# a_3125_n355#
+ a_1835_n355# a_n287_n300# a_n229_n355# a_n1061_n300# a_287_n355# a_n1003_n355# a_2809_n300#
+ a_745_n300# a_2093_n355# a_n3383_n300# a_n3325_n355# a_2551_n300# a_1319_n355#
X0 a_2809_n300# a_2609_n355# a_2551_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1 a_n2351_n300# a_n2551_n355# a_n2609_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X2 a_n2093_n300# a_n2293_n355# a_n2351_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3 a_n29_n300# a_n229_n355# a_n287_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X4 a_229_n300# a_29_n355# a_n29_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X5 a_3067_n300# a_2867_n355# a_2809_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 a_n1319_n300# a_n1519_n355# a_n1577_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_n545_n300# a_n745_n355# a_n803_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X8 a_2293_n300# a_2093_n355# a_2035_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X9 a_2551_n300# a_2351_n355# a_2293_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X10 a_n3125_n300# a_n3325_n355# a_n3383_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X11 a_n2867_n300# a_n3067_n355# a_n3125_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X12 a_n803_n300# a_n1003_n355# a_n1061_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_n287_n300# a_n487_n355# a_n545_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X14 a_n1577_n300# a_n1777_n355# a_n1835_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X15 a_1519_n300# a_1319_n355# a_1261_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 a_3325_n300# a_3125_n355# a_3067_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X17 a_n1061_n300# a_n1261_n355# a_n1319_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X18 a_745_n300# a_545_n355# a_487_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X19 a_1003_n300# a_803_n355# a_745_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X20 a_487_n300# a_287_n355# a_229_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X21 a_2035_n300# a_1835_n355# a_1777_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 a_n2609_n300# a_n2809_n355# a_n2867_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X23 a_1777_n300# a_1577_n355# a_1519_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_1261_n300# a_1061_n355# a_1003_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X25 a_n1835_n300# a_n2035_n355# a_n2093_n300# a_n3517_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
C0 a_n2093_n300# a_n2351_n300# 0.164742f
C1 a_n1061_n300# a_n803_n300# 0.164742f
C2 a_1777_n300# a_1519_n300# 0.164742f
C3 a_1519_n300# a_1261_n300# 0.164742f
C4 a_745_n300# a_487_n300# 0.164742f
C5 a_n287_n300# a_n29_n300# 0.164742f
C6 a_n287_n300# a_n545_n300# 0.164742f
C7 a_1777_n300# a_2035_n300# 0.164742f
C8 a_n2609_n300# a_n2351_n300# 0.164742f
C9 a_n2867_n300# a_n3125_n300# 0.164742f
C10 a_3325_n300# a_3067_n300# 0.164742f
C11 a_n1577_n300# a_n1319_n300# 0.164742f
C12 a_229_n300# a_n29_n300# 0.164742f
C13 a_n2867_n300# a_n2609_n300# 0.164742f
C14 a_487_n300# a_229_n300# 0.164742f
C15 a_1003_n300# a_1261_n300# 0.164742f
C16 a_n1835_n300# a_n2093_n300# 0.164742f
C17 a_2809_n300# a_2551_n300# 0.164742f
C18 a_n1835_n300# a_n1577_n300# 0.164742f
C19 a_n3125_n300# a_n3383_n300# 0.164742f
C20 a_745_n300# a_1003_n300# 0.164742f
C21 a_3067_n300# a_2809_n300# 0.164742f
C22 a_2293_n300# a_2551_n300# 0.164742f
C23 a_n545_n300# a_n803_n300# 0.164742f
C24 a_2293_n300# a_2035_n300# 0.164742f
C25 a_n1061_n300# a_n1319_n300# 0.164742f
C26 a_3325_n300# a_n3517_n522# 0.345442f
C27 a_3067_n300# a_n3517_n522# 0.111675f
C28 a_2809_n300# a_n3517_n522# 0.111675f
C29 a_2551_n300# a_n3517_n522# 0.111675f
C30 a_2293_n300# a_n3517_n522# 0.111675f
C31 a_2035_n300# a_n3517_n522# 0.111675f
C32 a_1777_n300# a_n3517_n522# 0.111675f
C33 a_1519_n300# a_n3517_n522# 0.111675f
C34 a_1261_n300# a_n3517_n522# 0.111675f
C35 a_1003_n300# a_n3517_n522# 0.111675f
C36 a_745_n300# a_n3517_n522# 0.111675f
C37 a_487_n300# a_n3517_n522# 0.111675f
C38 a_229_n300# a_n3517_n522# 0.111675f
C39 a_n29_n300# a_n3517_n522# 0.111675f
C40 a_n287_n300# a_n3517_n522# 0.111675f
C41 a_n545_n300# a_n3517_n522# 0.111675f
C42 a_n803_n300# a_n3517_n522# 0.111675f
C43 a_n1061_n300# a_n3517_n522# 0.111675f
C44 a_n1319_n300# a_n3517_n522# 0.111675f
C45 a_n1577_n300# a_n3517_n522# 0.111675f
C46 a_n1835_n300# a_n3517_n522# 0.111675f
C47 a_n2093_n300# a_n3517_n522# 0.111675f
C48 a_n2351_n300# a_n3517_n522# 0.111675f
C49 a_n2609_n300# a_n3517_n522# 0.111675f
C50 a_n2867_n300# a_n3517_n522# 0.111675f
C51 a_n3125_n300# a_n3517_n522# 0.111675f
C52 a_n3383_n300# a_n3517_n522# 0.345442f
C53 a_3125_n355# a_n3517_n522# 0.556766f
C54 a_2867_n355# a_n3517_n522# 0.502594f
C55 a_2609_n355# a_n3517_n522# 0.502594f
C56 a_2351_n355# a_n3517_n522# 0.502594f
C57 a_2093_n355# a_n3517_n522# 0.502594f
C58 a_1835_n355# a_n3517_n522# 0.502594f
C59 a_1577_n355# a_n3517_n522# 0.502594f
C60 a_1319_n355# a_n3517_n522# 0.502594f
C61 a_1061_n355# a_n3517_n522# 0.502594f
C62 a_803_n355# a_n3517_n522# 0.502594f
C63 a_545_n355# a_n3517_n522# 0.502594f
C64 a_287_n355# a_n3517_n522# 0.502594f
C65 a_29_n355# a_n3517_n522# 0.502594f
C66 a_n229_n355# a_n3517_n522# 0.502594f
C67 a_n487_n355# a_n3517_n522# 0.502594f
C68 a_n745_n355# a_n3517_n522# 0.502594f
C69 a_n1003_n355# a_n3517_n522# 0.502594f
C70 a_n1261_n355# a_n3517_n522# 0.502594f
C71 a_n1519_n355# a_n3517_n522# 0.502594f
C72 a_n1777_n355# a_n3517_n522# 0.502594f
C73 a_n2035_n355# a_n3517_n522# 0.502594f
C74 a_n2293_n355# a_n3517_n522# 0.502594f
C75 a_n2551_n355# a_n3517_n522# 0.502594f
C76 a_n2809_n355# a_n3517_n522# 0.502594f
C77 a_n3067_n355# a_n3517_n522# 0.502594f
C78 a_n3325_n355# a_n3517_n522# 0.556766f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2B7385 a_1261_n800# a_n1319_n800# a_1835_n855#
+ a_n287_n800# a_n229_n855# a_n1061_n800# a_287_n855# a_n1003_n855# a_2093_n855# a_745_n800#
+ a_1319_n855# a_1777_n800# a_n2293_n855# a_n2351_n800# a_1061_n855# a_229_n800# a_2035_n800#
+ a_n1577_n800# a_n1519_n855# a_n487_n855# a_n1261_n855# a_n545_n800# a_545_n855#
+ a_1003_n800# a_1577_n855# a_n2485_n1022# a_n29_n800# a_487_n800# a_2293_n800# a_29_n855#
+ a_n1777_n855# a_n1835_n800# a_n745_n855# a_n803_n800# a_1519_n800# a_n2093_n800#
+ a_803_n855# a_n2035_n855#
X0 a_n1577_n800# a_n1777_n855# a_n1835_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X1 a_1519_n800# a_1319_n855# a_1261_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2 a_n1061_n800# a_n1261_n855# a_n1319_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X3 a_1003_n800# a_803_n855# a_745_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X4 a_745_n800# a_545_n855# a_487_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X5 a_487_n800# a_287_n855# a_229_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X6 a_1777_n800# a_1577_n855# a_1519_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X7 a_2035_n800# a_1835_n855# a_1777_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X8 a_1261_n800# a_1061_n855# a_1003_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X9 a_n1835_n800# a_n2035_n855# a_n2093_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X10 a_n2093_n800# a_n2293_n855# a_n2351_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X11 a_n29_n800# a_n229_n855# a_n287_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X12 a_229_n800# a_29_n855# a_n29_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X13 a_n1319_n800# a_n1519_n855# a_n1577_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X14 a_n545_n800# a_n745_n855# a_n803_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X15 a_n287_n800# a_n487_n855# a_n545_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X16 a_2293_n800# a_2093_n855# a_2035_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X17 a_n803_n800# a_n1003_n855# a_n1061_n800# a_n2485_n1022# sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
C0 a_2093_n855# a_2035_n800# 0.176406f
C1 a_n287_n800# a_n487_n855# 0.176406f
C2 a_745_n800# a_803_n855# 0.176406f
C3 a_n1061_n800# a_n1319_n800# 0.437576f
C4 a_2293_n800# a_2035_n800# 0.437576f
C5 a_n2093_n800# a_n1835_n800# 0.437576f
C6 a_287_n855# a_229_n800# 0.176406f
C7 a_n1519_n855# a_n1577_n800# 0.176406f
C8 a_2293_n800# a_2093_n855# 0.176406f
C9 a_n29_n800# a_n229_n855# 0.176406f
C10 a_n2035_n855# a_n1835_n800# 0.176406f
C11 a_545_n855# a_487_n800# 0.176406f
C12 a_n1003_n855# a_n1061_n800# 0.176406f
C13 a_n2093_n800# a_n2035_n855# 0.176406f
C14 a_n745_n855# a_n803_n800# 0.176406f
C15 a_229_n800# a_n29_n800# 0.437576f
C16 a_n1577_n800# a_n1777_n855# 0.176406f
C17 a_745_n800# a_1003_n800# 0.437576f
C18 a_545_n855# a_745_n800# 0.176406f
C19 a_1835_n855# a_1777_n800# 0.176406f
C20 a_n1577_n800# a_n1319_n800# 0.437576f
C21 a_1777_n800# a_1519_n800# 0.437576f
C22 a_n2293_n855# a_n2351_n800# 0.176406f
C23 a_n29_n800# a_29_n855# 0.176406f
C24 a_229_n800# a_487_n800# 0.437576f
C25 a_n1777_n855# a_n1835_n800# 0.176406f
C26 a_n1261_n855# a_n1061_n800# 0.176406f
C27 a_1061_n855# a_1003_n800# 0.176406f
C28 a_1061_n855# a_1261_n800# 0.176406f
C29 a_1003_n800# a_803_n855# 0.176406f
C30 a_745_n800# a_487_n800# 0.437576f
C31 a_n803_n800# a_n1061_n800# 0.437576f
C32 a_n545_n800# a_n487_n855# 0.176406f
C33 a_1319_n855# a_1519_n800# 0.176406f
C34 a_1577_n855# a_1519_n800# 0.176406f
C35 a_1835_n855# a_2035_n800# 0.176406f
C36 a_1261_n800# a_1519_n800# 0.437576f
C37 a_n1261_n855# a_n1319_n800# 0.176406f
C38 a_1777_n800# a_1577_n855# 0.176406f
C39 a_n2293_n855# a_n2093_n800# 0.176406f
C40 a_n29_n800# a_n287_n800# 0.437576f
C41 a_1777_n800# a_2035_n800# 0.437576f
C42 a_n287_n800# a_n229_n855# 0.176406f
C43 a_229_n800# a_29_n855# 0.176406f
C44 a_n1577_n800# a_n1835_n800# 0.437576f
C45 a_n745_n855# a_n545_n800# 0.176406f
C46 a_n1519_n855# a_n1319_n800# 0.176406f
C47 a_1319_n855# a_1261_n800# 0.176406f
C48 a_n1003_n855# a_n803_n800# 0.176406f
C49 a_1261_n800# a_1003_n800# 0.437576f
C50 a_n545_n800# a_n803_n800# 0.437576f
C51 a_n2093_n800# a_n2351_n800# 0.437576f
C52 a_287_n855# a_487_n800# 0.176406f
C53 a_n545_n800# a_n287_n800# 0.437576f
C54 a_2293_n800# a_n2485_n1022# 0.86543f
C55 a_2035_n800# a_n2485_n1022# 0.248227f
C56 a_1777_n800# a_n2485_n1022# 0.248227f
C57 a_1519_n800# a_n2485_n1022# 0.248227f
C58 a_1261_n800# a_n2485_n1022# 0.248227f
C59 a_1003_n800# a_n2485_n1022# 0.248227f
C60 a_745_n800# a_n2485_n1022# 0.248227f
C61 a_487_n800# a_n2485_n1022# 0.248227f
C62 a_229_n800# a_n2485_n1022# 0.248227f
C63 a_n29_n800# a_n2485_n1022# 0.248227f
C64 a_n287_n800# a_n2485_n1022# 0.248227f
C65 a_n545_n800# a_n2485_n1022# 0.248227f
C66 a_n803_n800# a_n2485_n1022# 0.248227f
C67 a_n1061_n800# a_n2485_n1022# 0.248227f
C68 a_n1319_n800# a_n2485_n1022# 0.248227f
C69 a_n1577_n800# a_n2485_n1022# 0.248227f
C70 a_n1835_n800# a_n2485_n1022# 0.248227f
C71 a_n2093_n800# a_n2485_n1022# 0.248227f
C72 a_n2351_n800# a_n2485_n1022# 0.86543f
C73 a_2093_n855# a_n2485_n1022# 0.579228f
C74 a_1835_n855# a_n2485_n1022# 0.525056f
C75 a_1577_n855# a_n2485_n1022# 0.525056f
C76 a_1319_n855# a_n2485_n1022# 0.525056f
C77 a_1061_n855# a_n2485_n1022# 0.525056f
C78 a_803_n855# a_n2485_n1022# 0.525056f
C79 a_545_n855# a_n2485_n1022# 0.525056f
C80 a_287_n855# a_n2485_n1022# 0.525056f
C81 a_29_n855# a_n2485_n1022# 0.525056f
C82 a_n229_n855# a_n2485_n1022# 0.525056f
C83 a_n487_n855# a_n2485_n1022# 0.525056f
C84 a_n745_n855# a_n2485_n1022# 0.525056f
C85 a_n1003_n855# a_n2485_n1022# 0.525056f
C86 a_n1261_n855# a_n2485_n1022# 0.525056f
C87 a_n1519_n855# a_n2485_n1022# 0.525056f
C88 a_n1777_n855# a_n2485_n1022# 0.525056f
C89 a_n2035_n855# a_n2485_n1022# 0.525056f
C90 a_n2293_n855# a_n2485_n1022# 0.579228f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR a_n2093_n200# a_803_n255# a_n2035_n255#
+ a_n3841_n255# a_n5131_n255# a_1261_n200# a_n4357_n255# a_3583_n200# a_n1319_n200#
+ a_n4415_n200# a_4931_n255# a_3125_n255# a_1835_n255# a_n287_n200# a_n229_n255# a_4099_n200#
+ a_n1061_n200# a_287_n255# a_n1003_n255# a_2809_n200# a_745_n200# a_n3383_n200# a_2093_n255#
+ a_n3325_n255# a_2551_n200# a_3067_n200# a_4415_n255# a_1319_n255# a_4873_n200# a_1777_n200#
+ a_n2609_n200# a_n2293_n255# a_1061_n255# a_n5323_n422# a_n2351_n200# a_229_n200#
+ a_3383_n255# a_n1577_n200# a_n4673_n200# a_n1519_n255# a_n4615_n255# a_5131_n200#
+ a_3841_n200# a_2035_n200# a_n487_n255# a_n545_n200# a_n3899_n200# a_n5189_n200#
+ a_n1261_n255# a_4357_n200# a_2609_n255# a_545_n255# a_n3583_n255# a_n3641_n200#
+ a_2351_n255# a_1003_n200# a_n4099_n255# a_n4157_n200# a_4673_n255# a_1577_n255#
+ a_3325_n200# a_n2867_n200# a_n2809_n255# a_3899_n255# a_n2551_n255# a_487_n200#
+ a_n29_n200# a_n3067_n255# a_2293_n200# a_29_n255# a_n1777_n255# a_n4873_n255# a_n1835_n200#
+ a_n3125_n200# a_n4931_n200# a_3641_n255# a_4157_n255# a_n745_n255# a_n803_n200#
+ a_2867_n255# a_4615_n200# a_1519_n200#
X0 a_487_n200# a_287_n255# a_229_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_2035_n200# a_1835_n255# a_1777_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_4099_n200# a_3899_n255# a_3841_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n2609_n200# a_n2809_n255# a_n2867_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_1777_n200# a_1577_n255# a_1519_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_3841_n200# a_3641_n255# a_3583_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n4415_n200# a_n4615_n255# a_n4673_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_1261_n200# a_1061_n255# a_1003_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_3583_n200# a_3383_n255# a_3325_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n4157_n200# a_n4357_n255# a_n4415_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n3899_n200# a_n4099_n255# a_n4157_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1835_n200# a_n2035_n255# a_n2093_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_n4673_n200# a_n4873_n255# a_n4931_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_2809_n200# a_2609_n255# a_2551_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_n2351_n200# a_n2551_n255# a_n2609_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_4357_n200# a_4157_n255# a_4099_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_4615_n200# a_4415_n255# a_4357_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_n2093_n200# a_n2293_n255# a_n2351_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_n29_n200# a_n229_n255# a_n287_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_229_n200# a_29_n255# a_n29_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_3067_n200# a_2867_n255# a_2809_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X21 a_5131_n200# a_4931_n255# a_4873_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X22 a_4873_n200# a_4673_n255# a_4615_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X24 a_n545_n200# a_n745_n255# a_n803_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X25 a_2293_n200# a_2093_n255# a_2035_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 a_2551_n200# a_2351_n255# a_2293_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X27 a_n4931_n200# a_n5131_n255# a_n5189_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X28 a_n3125_n200# a_n3325_n255# a_n3383_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 a_n2867_n200# a_n3067_n255# a_n3125_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X31 a_n287_n200# a_n487_n255# a_n545_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X32 a_n3641_n200# a_n3841_n255# a_n3899_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_n1577_n200# a_n1777_n255# a_n1835_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 a_1519_n200# a_1319_n255# a_1261_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X35 a_n3383_n200# a_n3583_n255# a_n3641_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 a_3325_n200# a_3125_n255# a_3067_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X38 a_745_n200# a_545_n255# a_487_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X39 a_1003_n200# a_803_n255# a_745_n200# a_n5323_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
C0 a_487_n200# a_745_n200# 0.110175f
C1 a_3841_n200# a_4099_n200# 0.110175f
C2 a_1003_n200# a_745_n200# 0.110175f
C3 a_n545_n200# a_n287_n200# 0.110175f
C4 a_3325_n200# a_3583_n200# 0.110175f
C5 a_1003_n200# a_1261_n200# 0.110175f
C6 a_n3899_n200# a_n3641_n200# 0.110175f
C7 a_1519_n200# a_1777_n200# 0.110175f
C8 a_n803_n200# a_n545_n200# 0.110175f
C9 a_4873_n200# a_5131_n200# 0.110175f
C10 a_n4673_n200# a_n4931_n200# 0.110175f
C11 a_2551_n200# a_2809_n200# 0.110175f
C12 a_n29_n200# a_n287_n200# 0.110175f
C13 a_4099_n200# a_4357_n200# 0.110175f
C14 a_n2867_n200# a_n3125_n200# 0.110175f
C15 a_n1835_n200# a_n2093_n200# 0.110175f
C16 a_n1577_n200# a_n1319_n200# 0.110175f
C17 a_1777_n200# a_2035_n200# 0.110175f
C18 a_n3641_n200# a_n3383_n200# 0.110175f
C19 a_2551_n200# a_2293_n200# 0.110175f
C20 a_n4415_n200# a_n4673_n200# 0.110175f
C21 a_2809_n200# a_3067_n200# 0.110175f
C22 a_3583_n200# a_3841_n200# 0.110175f
C23 a_n5189_n200# a_n4931_n200# 0.110175f
C24 a_n3899_n200# a_n4157_n200# 0.110175f
C25 a_4357_n200# a_4615_n200# 0.110175f
C26 a_487_n200# a_229_n200# 0.110175f
C27 a_n1061_n200# a_n803_n200# 0.110175f
C28 a_n1061_n200# a_n1319_n200# 0.110175f
C29 a_n1577_n200# a_n1835_n200# 0.110175f
C30 a_2035_n200# a_2293_n200# 0.110175f
C31 a_n3125_n200# a_n3383_n200# 0.110175f
C32 a_3067_n200# a_3325_n200# 0.110175f
C33 a_1519_n200# a_1261_n200# 0.110175f
C34 a_n2351_n200# a_n2609_n200# 0.110175f
C35 a_229_n200# a_n29_n200# 0.110175f
C36 a_n2867_n200# a_n2609_n200# 0.110175f
C37 a_n4415_n200# a_n4157_n200# 0.110175f
C38 a_n2351_n200# a_n2093_n200# 0.110175f
C39 a_4615_n200# a_4873_n200# 0.110175f
C40 a_5131_n200# a_n5323_n422# 0.241444f
C41 a_n5189_n200# a_n5323_n422# 0.241444f
C42 a_4931_n255# a_n5323_n422# 0.55256f
C43 a_4673_n255# a_n5323_n422# 0.498389f
C44 a_4415_n255# a_n5323_n422# 0.498389f
C45 a_4157_n255# a_n5323_n422# 0.498389f
C46 a_3899_n255# a_n5323_n422# 0.498389f
C47 a_3641_n255# a_n5323_n422# 0.498389f
C48 a_3383_n255# a_n5323_n422# 0.498389f
C49 a_3125_n255# a_n5323_n422# 0.498389f
C50 a_2867_n255# a_n5323_n422# 0.498389f
C51 a_2609_n255# a_n5323_n422# 0.498389f
C52 a_2351_n255# a_n5323_n422# 0.498389f
C53 a_2093_n255# a_n5323_n422# 0.498389f
C54 a_1835_n255# a_n5323_n422# 0.498389f
C55 a_1577_n255# a_n5323_n422# 0.498389f
C56 a_1319_n255# a_n5323_n422# 0.498389f
C57 a_1061_n255# a_n5323_n422# 0.498389f
C58 a_803_n255# a_n5323_n422# 0.498389f
C59 a_545_n255# a_n5323_n422# 0.498389f
C60 a_287_n255# a_n5323_n422# 0.498389f
C61 a_29_n255# a_n5323_n422# 0.498389f
C62 a_n229_n255# a_n5323_n422# 0.498389f
C63 a_n487_n255# a_n5323_n422# 0.498389f
C64 a_n745_n255# a_n5323_n422# 0.498389f
C65 a_n1003_n255# a_n5323_n422# 0.498389f
C66 a_n1261_n255# a_n5323_n422# 0.498389f
C67 a_n1519_n255# a_n5323_n422# 0.498389f
C68 a_n1777_n255# a_n5323_n422# 0.498389f
C69 a_n2035_n255# a_n5323_n422# 0.498389f
C70 a_n2293_n255# a_n5323_n422# 0.498389f
C71 a_n2551_n255# a_n5323_n422# 0.498389f
C72 a_n2809_n255# a_n5323_n422# 0.498389f
C73 a_n3067_n255# a_n5323_n422# 0.498389f
C74 a_n3325_n255# a_n5323_n422# 0.498389f
C75 a_n3583_n255# a_n5323_n422# 0.498389f
C76 a_n3841_n255# a_n5323_n422# 0.498389f
C77 a_n4099_n255# a_n5323_n422# 0.498389f
C78 a_n4357_n255# a_n5323_n422# 0.498389f
C79 a_n4615_n255# a_n5323_n422# 0.498389f
C80 a_n4873_n255# a_n5323_n422# 0.498389f
C81 a_n5131_n255# a_n5323_n422# 0.55256f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_WK95DB a_n819_n450# a_n345_n450# a_29_n505# a_n129_n505#
+ a_187_n505# a_129_n450# a_n503_n450# a_n287_n505# a_345_n505# a_287_n450# a_n661_n450#
+ a_n445_n505# a_503_n505# a_445_n450# a_n603_n505# a_661_n505# a_603_n450# a_n761_n505#
+ a_761_n450# a_n953_n672# a_n29_n450# a_n187_n450#
X0 a_n345_n450# a_n445_n505# a_n503_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X1 a_129_n450# a_29_n505# a_n29_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X2 a_445_n450# a_345_n505# a_287_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X3 a_n503_n450# a_n603_n505# a_n661_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X4 a_n29_n450# a_n129_n505# a_n187_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X5 a_603_n450# a_503_n505# a_445_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X6 a_n661_n450# a_n761_n505# a_n819_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.5
X7 a_n187_n450# a_n287_n505# a_n345_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
X8 a_761_n450# a_661_n505# a_603_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.5
X9 a_287_n450# a_187_n505# a_129_n450# a_n953_n672# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.5
C0 a_n661_n450# a_n819_n450# 0.401603f
C1 a_n345_n450# a_n187_n450# 0.401603f
C2 a_445_n450# a_287_n450# 0.401603f
C3 a_n503_n450# a_n345_n450# 0.401603f
C4 a_n29_n450# a_129_n450# 0.401603f
C5 a_n29_n450# a_n187_n450# 0.401603f
C6 a_287_n450# a_129_n450# 0.401603f
C7 a_761_n450# a_603_n450# 0.401603f
C8 a_n503_n450# a_n661_n450# 0.401603f
C9 a_445_n450# a_603_n450# 0.401603f
C10 a_761_n450# a_n953_n672# 0.477209f
C11 a_603_n450# a_n953_n672# 0.104181f
C12 a_445_n450# a_n953_n672# 0.104181f
C13 a_287_n450# a_n953_n672# 0.104181f
C14 a_129_n450# a_n953_n672# 0.104181f
C15 a_n29_n450# a_n953_n672# 0.104181f
C16 a_n187_n450# a_n953_n672# 0.104181f
C17 a_n345_n450# a_n953_n672# 0.104181f
C18 a_n503_n450# a_n953_n672# 0.104181f
C19 a_n661_n450# a_n953_n672# 0.104181f
C20 a_n819_n450# a_n953_n672# 0.477209f
C21 a_661_n505# a_n953_n672# 0.334006f
C22 a_503_n505# a_n953_n672# 0.275258f
C23 a_345_n505# a_n953_n672# 0.275258f
C24 a_187_n505# a_n953_n672# 0.275258f
C25 a_29_n505# a_n953_n672# 0.275258f
C26 a_n129_n505# a_n953_n672# 0.275258f
C27 a_n287_n505# a_n953_n672# 0.275258f
C28 a_n445_n505# a_n953_n672# 0.275258f
C29 a_n603_n505# a_n953_n672# 0.275258f
C30 a_n761_n505# a_n953_n672# 0.334006f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3QL9S5 a_n50_n497# a_50_n400# w_n308_n697# a_n108_n400#
X0 a_50_n400# a_n50_n497# a_n108_n400# w_n308_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
C0 a_50_n400# w_n308_n697# 0.249352f
C1 a_n108_n400# w_n308_n697# 0.249352f
C2 a_n50_n497# w_n308_n697# 0.280349f
C3 a_n108_n400# a_50_n400# 0.357178f
C4 a_50_n400# 0 0.180042f
C5 a_n108_n400# 0 0.180042f
C6 a_n50_n497# 0 0.168405f
C7 w_n308_n697# 0 3.39795f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PGZBW9 a_1061_n655# a_n2293_n655# a_n2351_n600#
+ a_229_n600# a_n1577_n600# a_n1519_n655# a_2035_n600# a_n487_n655# a_n1261_n655#
+ a_n545_n600# a_2609_n655# a_545_n655# a_2351_n655# a_n3517_n822# a_1003_n600# a_1577_n655#
+ a_n2867_n600# a_n2809_n655# a_3325_n600# a_n2551_n655# a_n29_n600# a_487_n600# a_n1777_n655#
+ a_n3067_n655# a_2293_n600# a_n3125_n600# a_29_n655# a_n1835_n600# a_2867_n655# a_n745_n655#
+ a_n803_n600# a_1519_n600# a_n2093_n600# a_803_n655# a_n2035_n655# a_1261_n600# a_3125_n655#
+ a_n1319_n600# a_1835_n655# a_n287_n600# a_n1061_n600# a_n229_n655# a_n1003_n655#
+ a_287_n655# a_2809_n600# a_2093_n655# a_745_n600# a_n3383_n600# a_n3325_n655# a_2551_n600#
+ a_3067_n600# a_1777_n600# a_n2609_n600# a_1319_n655#
X0 a_2809_n600# a_2609_n655# a_2551_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n655# a_n2609_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n655# a_n2351_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_229_n600# a_29_n655# a_n29_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_n29_n600# a_n229_n655# a_n287_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n655# a_2809_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n655# a_n1577_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n655# a_2293_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n655# a_n3383_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X9 a_n545_n600# a_n745_n655# a_n803_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n655# a_n545_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n655# a_2035_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n655# a_n3125_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n655# a_n1061_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n1577_n600# a_n1777_n655# a_n1835_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X15 a_1519_n600# a_1319_n655# a_1261_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_n1061_n600# a_n1261_n655# a_n1319_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_3325_n600# a_3125_n655# a_3067_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X18 a_1003_n600# a_803_n655# a_745_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_745_n600# a_545_n655# a_487_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_487_n600# a_287_n655# a_229_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_2035_n600# a_1835_n655# a_1777_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_n2609_n600# a_n2809_n655# a_n2867_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_1777_n600# a_1577_n655# a_1519_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1261_n600# a_1061_n655# a_1003_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_n1835_n600# a_n2035_n655# a_n2093_n600# a_n3517_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
C0 a_3125_n655# a_3325_n600# 0.133664f
C1 a_n2809_n655# a_n2867_n600# 0.133664f
C2 a_n1519_n655# a_n1319_n600# 0.133664f
C3 a_2093_n655# a_2035_n600# 0.133664f
C4 a_2293_n600# a_2035_n600# 0.328443f
C5 a_n2351_n600# a_n2609_n600# 0.328443f
C6 a_1777_n600# a_2035_n600# 0.328443f
C7 a_1777_n600# a_1835_n655# 0.133664f
C8 a_803_n655# a_1003_n600# 0.133664f
C9 a_n2293_n655# a_n2351_n600# 0.133664f
C10 a_1519_n600# a_1319_n655# 0.133664f
C11 a_n1835_n600# a_n2035_n655# 0.133664f
C12 a_n2093_n600# a_n2035_n655# 0.133664f
C13 a_n1577_n600# a_n1777_n655# 0.133664f
C14 a_n2809_n655# a_n2609_n600# 0.133664f
C15 a_745_n600# a_1003_n600# 0.328443f
C16 a_229_n600# a_487_n600# 0.328443f
C17 a_n3067_n655# a_n2867_n600# 0.133664f
C18 a_2035_n600# a_1835_n655# 0.133664f
C19 a_n287_n600# a_n29_n600# 0.328443f
C20 a_n3325_n655# a_n3125_n600# 0.133664f
C21 a_229_n600# a_n29_n600# 0.328443f
C22 a_2551_n600# a_2609_n655# 0.133664f
C23 a_n1577_n600# a_n1835_n600# 0.328443f
C24 a_n229_n655# a_n29_n600# 0.133664f
C25 a_1061_n655# a_1003_n600# 0.133664f
C26 a_29_n655# a_n29_n600# 0.133664f
C27 a_1577_n655# a_1777_n600# 0.133664f
C28 a_n2351_n600# a_n2093_n600# 0.328443f
C29 a_n803_n600# a_n745_n655# 0.133664f
C30 a_n3383_n600# a_n3325_n655# 0.133664f
C31 a_n2293_n655# a_n2093_n600# 0.133664f
C32 a_2867_n655# a_2809_n600# 0.133664f
C33 a_3067_n600# a_2809_n600# 0.328443f
C34 a_3067_n600# a_2867_n655# 0.133664f
C35 a_n1777_n655# a_n1835_n600# 0.133664f
C36 a_n487_n655# a_n545_n600# 0.133664f
C37 a_n487_n655# a_n287_n600# 0.133664f
C38 a_n1577_n600# a_n1319_n600# 0.328443f
C39 a_n1577_n600# a_n1519_n655# 0.133664f
C40 a_n545_n600# a_n745_n655# 0.133664f
C41 a_n3383_n600# a_n3125_n600# 0.328443f
C42 a_545_n655# a_487_n600# 0.133664f
C43 a_1319_n655# a_1261_n600# 0.133664f
C44 a_1519_n600# a_1777_n600# 0.328443f
C45 a_n803_n600# a_n545_n600# 0.328443f
C46 a_n1061_n600# a_n803_n600# 0.328443f
C47 a_229_n600# a_287_n655# 0.133664f
C48 a_n2093_n600# a_n1835_n600# 0.328443f
C49 a_n2867_n600# a_n3125_n600# 0.328443f
C50 a_1061_n655# a_1261_n600# 0.133664f
C51 a_1519_n600# a_1261_n600# 0.328443f
C52 a_n1261_n655# a_n1061_n600# 0.133664f
C53 a_n1003_n655# a_n803_n600# 0.133664f
C54 a_2551_n600# a_2809_n600# 0.328443f
C55 a_745_n600# a_487_n600# 0.328443f
C56 a_n287_n600# a_n545_n600# 0.328443f
C57 a_1261_n600# a_1003_n600# 0.328443f
C58 a_3067_n600# a_3325_n600# 0.328443f
C59 a_545_n655# a_745_n600# 0.133664f
C60 a_n2351_n600# a_n2551_n655# 0.133664f
C61 a_2351_n655# a_2293_n600# 0.133664f
C62 a_3125_n655# a_3067_n600# 0.133664f
C63 a_n1261_n655# a_n1319_n600# 0.133664f
C64 a_n229_n655# a_n287_n600# 0.133664f
C65 a_n2551_n655# a_n2609_n600# 0.133664f
C66 a_2551_n600# a_2351_n655# 0.133664f
C67 a_745_n600# a_803_n655# 0.133664f
C68 a_n1003_n655# a_n1061_n600# 0.133664f
C69 a_229_n600# a_29_n655# 0.133664f
C70 a_n1061_n600# a_n1319_n600# 0.328443f
C71 a_2093_n655# a_2293_n600# 0.133664f
C72 a_287_n655# a_487_n600# 0.133664f
C73 a_1577_n655# a_1519_n600# 0.133664f
C74 a_2551_n600# a_2293_n600# 0.328443f
C75 a_n2867_n600# a_n2609_n600# 0.328443f
C76 a_n3067_n655# a_n3125_n600# 0.133664f
C77 a_2609_n655# a_2809_n600# 0.133664f
C78 a_3325_n600# a_n3517_n822# 0.657435f
C79 a_3067_n600# a_n3517_n822# 0.193606f
C80 a_2809_n600# a_n3517_n822# 0.193606f
C81 a_2551_n600# a_n3517_n822# 0.193606f
C82 a_2293_n600# a_n3517_n822# 0.193606f
C83 a_2035_n600# a_n3517_n822# 0.193606f
C84 a_1777_n600# a_n3517_n822# 0.193606f
C85 a_1519_n600# a_n3517_n822# 0.193606f
C86 a_1261_n600# a_n3517_n822# 0.193606f
C87 a_1003_n600# a_n3517_n822# 0.193606f
C88 a_745_n600# a_n3517_n822# 0.193606f
C89 a_487_n600# a_n3517_n822# 0.193606f
C90 a_229_n600# a_n3517_n822# 0.193606f
C91 a_n29_n600# a_n3517_n822# 0.193606f
C92 a_n287_n600# a_n3517_n822# 0.193606f
C93 a_n545_n600# a_n3517_n822# 0.193606f
C94 a_n803_n600# a_n3517_n822# 0.193606f
C95 a_n1061_n600# a_n3517_n822# 0.193606f
C96 a_n1319_n600# a_n3517_n822# 0.193606f
C97 a_n1577_n600# a_n3517_n822# 0.193606f
C98 a_n1835_n600# a_n3517_n822# 0.193606f
C99 a_n2093_n600# a_n3517_n822# 0.193606f
C100 a_n2351_n600# a_n3517_n822# 0.193606f
C101 a_n2609_n600# a_n3517_n822# 0.193606f
C102 a_n2867_n600# a_n3517_n822# 0.193606f
C103 a_n3125_n600# a_n3517_n822# 0.193606f
C104 a_n3383_n600# a_n3517_n822# 0.657435f
C105 a_3125_n655# a_n3517_n822# 0.562598f
C106 a_2867_n655# a_n3517_n822# 0.508426f
C107 a_2609_n655# a_n3517_n822# 0.508426f
C108 a_2351_n655# a_n3517_n822# 0.508426f
C109 a_2093_n655# a_n3517_n822# 0.508426f
C110 a_1835_n655# a_n3517_n822# 0.508426f
C111 a_1577_n655# a_n3517_n822# 0.508426f
C112 a_1319_n655# a_n3517_n822# 0.508426f
C113 a_1061_n655# a_n3517_n822# 0.508426f
C114 a_803_n655# a_n3517_n822# 0.508426f
C115 a_545_n655# a_n3517_n822# 0.508426f
C116 a_287_n655# a_n3517_n822# 0.508426f
C117 a_29_n655# a_n3517_n822# 0.508426f
C118 a_n229_n655# a_n3517_n822# 0.508426f
C119 a_n487_n655# a_n3517_n822# 0.508426f
C120 a_n745_n655# a_n3517_n822# 0.508426f
C121 a_n1003_n655# a_n3517_n822# 0.508426f
C122 a_n1261_n655# a_n3517_n822# 0.508426f
C123 a_n1519_n655# a_n3517_n822# 0.508426f
C124 a_n1777_n655# a_n3517_n822# 0.508426f
C125 a_n2035_n655# a_n3517_n822# 0.508426f
C126 a_n2293_n655# a_n3517_n822# 0.508426f
C127 a_n2551_n655# a_n3517_n822# 0.508426f
C128 a_n2809_n655# a_n3517_n822# 0.508426f
C129 a_n3067_n655# a_n3517_n822# 0.508426f
C130 a_n3325_n655# a_n3517_n822# 0.562598f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD a_761_n400# a_503_n464# a_n29_n400# a_n603_n464#
+ a_661_n464# a_n187_n400# a_n761_n464# a_n819_n400# a_n345_n400# a_129_n400# a_n503_n400#
+ w_n1019_n697# a_287_n400# a_n661_n400# a_29_n464# a_n129_n464# a_187_n464# a_445_n400#
+ a_n287_n464# a_345_n464# a_603_n400# a_n445_n464#
X0 a_n503_n400# a_n603_n464# a_n661_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X1 a_n29_n400# a_n129_n464# a_n187_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X2 a_603_n400# a_503_n464# a_445_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X3 a_n661_n400# a_n761_n464# a_n819_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X4 a_n187_n400# a_n287_n464# a_n345_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X5 a_761_n400# a_661_n464# a_603_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X6 a_287_n400# a_187_n464# a_129_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X7 a_n345_n400# a_n445_n464# a_n503_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X8 a_129_n400# a_29_n464# a_n29_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
X9 a_445_n400# a_345_n464# a_287_n400# w_n1019_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=0.5
C0 a_n129_n464# w_n1019_n697# 0.180946f
C1 a_503_n464# w_n1019_n697# 0.180946f
C2 a_129_n400# a_n29_n400# 0.357178f
C3 w_n1019_n697# a_187_n464# 0.180946f
C4 a_661_n464# w_n1019_n697# 0.220136f
C5 a_n345_n400# a_n503_n400# 0.357178f
C6 a_129_n400# a_287_n400# 0.357178f
C7 a_603_n400# a_761_n400# 0.357178f
C8 a_445_n400# a_603_n400# 0.357178f
C9 a_n187_n400# a_n29_n400# 0.357178f
C10 a_n503_n400# a_n661_n400# 0.357178f
C11 w_n1019_n697# a_n603_n464# 0.180946f
C12 w_n1019_n697# a_n819_n400# 0.249352f
C13 a_n187_n400# a_n345_n400# 0.357178f
C14 a_n445_n464# w_n1019_n697# 0.180946f
C15 a_n661_n400# a_n819_n400# 0.357178f
C16 w_n1019_n697# a_761_n400# 0.249352f
C17 a_345_n464# w_n1019_n697# 0.180946f
C18 a_445_n400# a_287_n400# 0.357178f
C19 w_n1019_n697# a_29_n464# 0.180946f
C20 w_n1019_n697# a_n287_n464# 0.180946f
C21 a_n761_n464# w_n1019_n697# 0.220136f
C22 a_761_n400# 0 0.180042f
C23 a_n819_n400# 0 0.180042f
C24 a_661_n464# 0 0.125675f
C25 a_503_n464# 0 0.102602f
C26 a_345_n464# 0 0.102602f
C27 a_187_n464# 0 0.102602f
C28 a_29_n464# 0 0.102602f
C29 a_n129_n464# 0 0.102602f
C30 a_n287_n464# 0 0.102602f
C31 a_n445_n464# 0 0.102602f
C32 a_n603_n464# 0 0.102602f
C33 a_n761_n464# 0 0.125675f
C34 w_n1019_n697# 0 10.2323f
.ends

.subckt sky130_fd_pr__res_generic_po_U7N8A7 a_n719_n1060# a_n589_n930# a_n467_n930#
+ a_n345_n930# a_265_500# a_n223_n930# a_n101_n930# a_n223_500# a_21_500# a_n467_500#
+ a_509_500# a_143_500# a_509_n930# a_387_n930# a_387_500# a_265_n930# a_n101_500#
+ a_143_n930# a_n345_500# a_n589_500# a_21_n930#
R0 a_265_500# a_265_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R1 a_509_500# a_509_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R2 a_n467_500# a_n467_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R3 a_n101_500# a_n101_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R4 a_21_500# a_21_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R5 a_143_500# a_143_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R6 a_n345_500# a_n345_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R7 a_387_500# a_387_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R8 a_n589_500# a_n589_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
R9 a_n223_500# a_n223_n930# sky130_fd_pr__res_generic_po w=0.4 l=5
C0 a_n101_n930# a_n223_n930# 0.438212f
C1 a_265_n930# a_143_n930# 0.438212f
C2 a_387_500# a_509_500# 0.438212f
C3 a_n345_500# a_n467_500# 0.438212f
C4 a_21_n930# a_n101_n930# 0.438212f
C5 a_n223_500# a_n101_500# 0.438212f
C6 a_265_500# a_143_500# 0.438212f
C7 a_n345_500# a_n223_500# 0.438212f
C8 a_n345_n930# a_n467_n930# 0.438212f
C9 a_509_n930# a_387_n930# 0.438212f
C10 a_265_n930# a_387_n930# 0.438212f
C11 a_21_n930# a_143_n930# 0.438212f
C12 a_n467_500# a_n589_500# 0.438212f
C13 a_21_500# a_n101_500# 0.438212f
C14 a_387_500# a_265_500# 0.438212f
C15 a_21_500# a_143_500# 0.438212f
C16 a_n467_n930# a_n589_n930# 0.438212f
C17 a_n345_n930# a_n223_n930# 0.438212f
C18 a_509_n930# a_n719_n1060# 0.535751f
C19 a_509_500# a_n719_n1060# 0.535751f
C20 a_387_n930# a_n719_n1060# 0.280864f
C21 a_387_500# a_n719_n1060# 0.280864f
C22 a_265_n930# a_n719_n1060# 0.280864f
C23 a_265_500# a_n719_n1060# 0.280864f
C24 a_143_n930# a_n719_n1060# 0.280864f
C25 a_143_500# a_n719_n1060# 0.280864f
C26 a_21_n930# a_n719_n1060# 0.280864f
C27 a_21_500# a_n719_n1060# 0.280864f
C28 a_n101_n930# a_n719_n1060# 0.280864f
C29 a_n101_500# a_n719_n1060# 0.280864f
C30 a_n223_n930# a_n719_n1060# 0.280864f
C31 a_n223_500# a_n719_n1060# 0.280864f
C32 a_n345_n930# a_n719_n1060# 0.280864f
C33 a_n345_500# a_n719_n1060# 0.280864f
C34 a_n467_n930# a_n719_n1060# 0.280864f
C35 a_n467_500# a_n719_n1060# 0.280864f
C36 a_n589_n930# a_n719_n1060# 0.535751f
C37 a_n589_500# a_n719_n1060# 0.535751f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QSKB8C a_287_n464# a_n1003_n464# a_n2867_n400#
+ a_n4157_n400# a_2093_n464# a_3325_n400# a_n3325_n464# a_487_n400# a_n29_n400# a_4415_n464#
+ a_1319_n464# a_2293_n400# a_n1835_n400# a_n3125_n400# a_n2293_n464# a_n4931_n400#
+ a_1061_n464# a_1519_n400# a_n803_n400# a_3383_n464# a_4615_n400# a_n2093_n400# a_n1519_n464#
+ a_n4615_n464# a_1261_n400# a_n487_n464# a_n1261_n464# w_n5131_n697# a_n1319_n400#
+ a_2609_n464# a_545_n464# a_3583_n400# a_n287_n400# a_n4415_n400# a_n3583_n464# a_4099_n400#
+ a_n1061_n400# a_2351_n464# a_n4099_n464# a_2809_n400# a_4673_n464# a_1577_n464#
+ a_745_n400# a_n3383_n400# a_n2809_n464# a_2551_n400# a_3899_n464# a_n2551_n464#
+ a_4873_n400# a_3067_n400# a_1777_n400# a_n2609_n400# a_n3067_n464# a_3641_n464#
+ a_29_n464# a_n1777_n464# a_n4873_n464# a_n2351_n400# a_4157_n464# a_n745_n464# a_229_n400#
+ a_n1577_n400# a_n4673_n400# a_2867_n464# a_2035_n400# a_803_n464# a_n2035_n464#
+ a_3841_n400# a_n3841_n464# a_4357_n400# a_n545_n400# a_n3899_n400# a_3125_n464#
+ a_n4357_n464# a_1835_n464# a_1003_n400# a_n3641_n400# a_n229_n464#
X0 a_3067_n400# a_2867_n464# a_2809_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_4873_n400# a_4673_n464# a_4615_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_n545_n400# a_n745_n464# a_n803_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_2293_n400# a_2093_n464# a_2035_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_2551_n400# a_2351_n464# a_2293_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n3125_n400# a_n3325_n464# a_n3383_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n2867_n400# a_n3067_n464# a_n3125_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_n287_n400# a_n487_n464# a_n545_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n3641_n400# a_n3841_n464# a_n3899_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_n1577_n400# a_n1777_n464# a_n1835_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_1519_n400# a_1319_n464# a_1261_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_n3383_n400# a_n3583_n464# a_n3641_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_3325_n400# a_3125_n464# a_3067_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_1003_n400# a_803_n464# a_745_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_487_n400# a_287_n464# a_229_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_745_n400# a_545_n464# a_487_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_2035_n400# a_1835_n464# a_1777_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_4099_n400# a_3899_n464# a_3841_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_n2609_n400# a_n2809_n464# a_n2867_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X22 a_1777_n400# a_1577_n464# a_1519_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X23 a_3841_n400# a_3641_n464# a_3583_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X24 a_n4415_n400# a_n4615_n464# a_n4673_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 a_1261_n400# a_1061_n464# a_1003_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X26 a_3583_n400# a_3383_n464# a_3325_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X27 a_n4157_n400# a_n4357_n464# a_n4415_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X28 a_n3899_n400# a_n4099_n464# a_n4157_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X29 a_n1835_n400# a_n2035_n464# a_n2093_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X30 a_n4673_n400# a_n4873_n464# a_n4931_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X31 a_2809_n400# a_2609_n464# a_2551_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X32 a_n2351_n400# a_n2551_n464# a_n2609_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X33 a_4357_n400# a_4157_n464# a_4099_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X34 a_4615_n400# a_4415_n464# a_4357_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X35 a_n2093_n400# a_n2293_n464# a_n2351_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X36 a_n29_n400# a_n229_n464# a_n287_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X37 a_229_n400# a_29_n464# a_n29_n400# w_n5131_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
C0 a_3325_n400# a_3583_n400# 0.219309f
C1 a_487_n400# a_745_n400# 0.219309f
C2 w_n5131_n697# a_n2293_n464# 0.307639f
C3 a_3067_n400# a_3325_n400# 0.219309f
C4 w_n5131_n697# a_2351_n464# 0.307639f
C5 a_n1319_n400# a_n1061_n400# 0.219309f
C6 w_n5131_n697# a_n1519_n464# 0.307639f
C7 a_2809_n400# a_3067_n400# 0.219309f
C8 a_1519_n400# a_1777_n400# 0.219309f
C9 w_n5131_n697# a_29_n464# 0.307639f
C10 w_n5131_n697# a_n229_n464# 0.307639f
C11 a_2035_n400# a_1777_n400# 0.219309f
C12 a_n3899_n400# a_n4157_n400# 0.219309f
C13 w_n5131_n697# a_n1777_n464# 0.307639f
C14 w_n5131_n697# a_2867_n464# 0.307639f
C15 w_n5131_n697# a_1835_n464# 0.307639f
C16 a_2035_n400# a_2293_n400# 0.219309f
C17 a_n3125_n400# a_n2867_n400# 0.219309f
C18 a_4357_n400# a_4615_n400# 0.219309f
C19 a_545_n464# w_n5131_n697# 0.307639f
C20 w_n5131_n697# a_n3325_n464# 0.307639f
C21 a_487_n400# a_229_n400# 0.219309f
C22 w_n5131_n697# a_4673_n464# 0.34286f
C23 a_3583_n400# a_3841_n400# 0.219309f
C24 a_n545_n400# a_n287_n400# 0.219309f
C25 a_n2035_n464# w_n5131_n697# 0.307639f
C26 w_n5131_n697# a_n745_n464# 0.307639f
C27 a_n2093_n400# a_n2351_n400# 0.219309f
C28 a_n4157_n400# a_n4415_n400# 0.219309f
C29 w_n5131_n697# a_n4357_n464# 0.307639f
C30 w_n5131_n697# a_n2551_n464# 0.307639f
C31 w_n5131_n697# a_n4615_n464# 0.307639f
C32 w_n5131_n697# a_3641_n464# 0.307639f
C33 a_n3583_n464# w_n5131_n697# 0.307639f
C34 a_2293_n400# a_2551_n400# 0.219309f
C35 a_1003_n400# a_1261_n400# 0.219309f
C36 a_745_n400# a_1003_n400# 0.219309f
C37 w_n5131_n697# a_2609_n464# 0.307639f
C38 w_n5131_n697# a_n1261_n464# 0.307639f
C39 w_n5131_n697# a_287_n464# 0.307639f
C40 a_n545_n400# a_n803_n400# 0.219309f
C41 a_4615_n400# a_4873_n400# 0.219309f
C42 w_n5131_n697# a_803_n464# 0.307639f
C43 w_n5131_n697# a_n2809_n464# 0.307639f
C44 a_n2609_n400# a_n2351_n400# 0.219309f
C45 a_n2867_n400# a_n2609_n400# 0.219309f
C46 a_n29_n400# a_n287_n400# 0.219309f
C47 a_n29_n400# a_229_n400# 0.219309f
C48 a_n4673_n400# a_n4931_n400# 0.219309f
C49 a_3841_n400# a_4099_n400# 0.219309f
C50 w_n5131_n697# a_n487_n464# 0.307639f
C51 a_n3899_n400# a_n3641_n400# 0.219309f
C52 w_n5131_n697# a_2093_n464# 0.307639f
C53 a_n4099_n464# w_n5131_n697# 0.307639f
C54 w_n5131_n697# a_n3841_n464# 0.307639f
C55 a_n1319_n400# a_n1577_n400# 0.219309f
C56 w_n5131_n697# a_3383_n464# 0.307639f
C57 w_n5131_n697# a_4157_n464# 0.307639f
C58 w_n5131_n697# a_1577_n464# 0.307639f
C59 w_n5131_n697# a_n4873_n464# 0.34286f
C60 a_2551_n400# a_2809_n400# 0.219309f
C61 a_1261_n400# a_1519_n400# 0.219309f
C62 w_n5131_n697# a_1061_n464# 0.307639f
C63 w_n5131_n697# a_4415_n464# 0.307639f
C64 a_n2093_n400# a_n1835_n400# 0.219309f
C65 w_n5131_n697# a_n3067_n464# 0.307639f
C66 w_n5131_n697# a_n1003_n464# 0.307639f
C67 w_n5131_n697# a_4873_n400# 0.249341f
C68 w_n5131_n697# a_3899_n464# 0.307639f
C69 w_n5131_n697# a_1319_n464# 0.307639f
C70 w_n5131_n697# a_3125_n464# 0.307639f
C71 a_n3125_n400# a_n3383_n400# 0.219309f
C72 a_4099_n400# a_4357_n400# 0.219309f
C73 a_n3383_n400# a_n3641_n400# 0.219309f
C74 a_n4673_n400# a_n4415_n400# 0.219309f
C75 a_n803_n400# a_n1061_n400# 0.219309f
C76 w_n5131_n697# a_n4931_n400# 0.249341f
C77 a_n1577_n400# a_n1835_n400# 0.219309f
C78 a_4873_n400# 0 0.201515f
C79 a_4615_n400# 0 0.116864f
C80 a_4357_n400# 0 0.116864f
C81 a_4099_n400# 0 0.116864f
C82 a_3841_n400# 0 0.116864f
C83 a_3583_n400# 0 0.116864f
C84 a_3325_n400# 0 0.116864f
C85 a_3067_n400# 0 0.116864f
C86 a_2809_n400# 0 0.116864f
C87 a_2551_n400# 0 0.116864f
C88 a_2293_n400# 0 0.116864f
C89 a_2035_n400# 0 0.116864f
C90 a_1777_n400# 0 0.116864f
C91 a_1519_n400# 0 0.116864f
C92 a_1261_n400# 0 0.116864f
C93 a_1003_n400# 0 0.116864f
C94 a_745_n400# 0 0.116864f
C95 a_487_n400# 0 0.116864f
C96 a_229_n400# 0 0.116864f
C97 a_n29_n400# 0 0.116864f
C98 a_n287_n400# 0 0.116864f
C99 a_n545_n400# 0 0.116864f
C100 a_n803_n400# 0 0.116864f
C101 a_n1061_n400# 0 0.116864f
C102 a_n1319_n400# 0 0.116864f
C103 a_n1577_n400# 0 0.116864f
C104 a_n1835_n400# 0 0.116864f
C105 a_n2093_n400# 0 0.116864f
C106 a_n2351_n400# 0 0.116864f
C107 a_n2609_n400# 0 0.116864f
C108 a_n2867_n400# 0 0.116864f
C109 a_n3125_n400# 0 0.116864f
C110 a_n3383_n400# 0 0.116864f
C111 a_n3641_n400# 0 0.116864f
C112 a_n3899_n400# 0 0.116864f
C113 a_n4157_n400# 0 0.116864f
C114 a_n4415_n400# 0 0.116864f
C115 a_n4673_n400# 0 0.116864f
C116 a_n4931_n400# 0 0.201515f
C117 a_4673_n464# 0 0.233871f
C118 a_4415_n464# 0 0.211442f
C119 a_4157_n464# 0 0.211442f
C120 a_3899_n464# 0 0.211442f
C121 a_3641_n464# 0 0.211442f
C122 a_3383_n464# 0 0.211442f
C123 a_3125_n464# 0 0.211442f
C124 a_2867_n464# 0 0.211442f
C125 a_2609_n464# 0 0.211442f
C126 a_2351_n464# 0 0.211442f
C127 a_2093_n464# 0 0.211442f
C128 a_1835_n464# 0 0.211442f
C129 a_1577_n464# 0 0.211442f
C130 a_1319_n464# 0 0.211442f
C131 a_1061_n464# 0 0.211442f
C132 a_803_n464# 0 0.211442f
C133 a_545_n464# 0 0.211442f
C134 a_287_n464# 0 0.211442f
C135 a_29_n464# 0 0.211442f
C136 a_n229_n464# 0 0.211442f
C137 a_n487_n464# 0 0.211442f
C138 a_n745_n464# 0 0.211442f
C139 a_n1003_n464# 0 0.211442f
C140 a_n1261_n464# 0 0.211442f
C141 a_n1519_n464# 0 0.211442f
C142 a_n1777_n464# 0 0.211442f
C143 a_n2035_n464# 0 0.211442f
C144 a_n2293_n464# 0 0.211442f
C145 a_n2551_n464# 0 0.211442f
C146 a_n2809_n464# 0 0.211442f
C147 a_n3067_n464# 0 0.211442f
C148 a_n3325_n464# 0 0.211442f
C149 a_n3583_n464# 0 0.211442f
C150 a_n3841_n464# 0 0.211442f
C151 a_n4099_n464# 0 0.211442f
C152 a_n4357_n464# 0 0.211442f
C153 a_n4615_n464# 0 0.211442f
C154 a_n4873_n464# 0 0.233871f
C155 w_n5131_n697# 0 49.563602f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_QRKB8C a_287_n464# a_n1003_n464# a_n2867_n400#
+ a_n4157_n400# a_2093_n464# a_3325_n400# a_n3325_n464# a_487_n400# a_n29_n400# a_4415_n464#
+ a_1319_n464# a_2293_n400# a_n1835_n400# a_n3125_n400# a_n2293_n464# a_1061_n464#
+ w_n4873_n697# a_1519_n400# a_n803_n400# a_3383_n464# a_4615_n400# a_n2093_n400#
+ a_n1519_n464# a_n4615_n464# a_1261_n400# a_n487_n464# a_n1261_n464# a_n1319_n400#
+ a_2609_n464# a_545_n464# a_3583_n400# a_n287_n400# a_n4415_n400# a_n3583_n464# a_4099_n400#
+ a_n1061_n400# a_2351_n464# a_n4099_n464# a_2809_n400# a_1577_n464# a_745_n400# a_n3383_n400#
+ a_n2809_n464# a_2551_n400# a_3899_n464# a_n2551_n464# a_3067_n400# a_1777_n400#
+ a_n2609_n400# a_n3067_n464# a_3641_n464# a_29_n464# a_n1777_n464# a_n2351_n400#
+ a_4157_n464# a_n745_n464# a_229_n400# a_n1577_n400# a_n4673_n400# a_2867_n464# a_2035_n400#
+ a_803_n464# a_n2035_n464# a_3841_n400# a_n3841_n464# a_4357_n400# a_n545_n400# a_n3899_n400#
+ a_3125_n464# a_n4357_n464# a_1835_n464# a_1003_n400# a_n3641_n400# a_n229_n464#
X0 a_3067_n400# a_2867_n464# a_2809_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X1 a_n1319_n400# a_n1519_n464# a_n1577_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2 a_n545_n400# a_n745_n464# a_n803_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X3 a_2293_n400# a_2093_n464# a_2035_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X4 a_2551_n400# a_2351_n464# a_2293_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X5 a_n3125_n400# a_n3325_n464# a_n3383_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X6 a_n2867_n400# a_n3067_n464# a_n3125_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X7 a_n803_n400# a_n1003_n464# a_n1061_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X8 a_n287_n400# a_n487_n464# a_n545_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X9 a_n3641_n400# a_n3841_n464# a_n3899_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X10 a_n1577_n400# a_n1777_n464# a_n1835_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X11 a_1519_n400# a_1319_n464# a_1261_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X12 a_n3383_n400# a_n3583_n464# a_n3641_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X13 a_3325_n400# a_3125_n464# a_3067_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X14 a_n1061_n400# a_n1261_n464# a_n1319_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X15 a_1003_n400# a_803_n464# a_745_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X16 a_487_n400# a_287_n464# a_229_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X17 a_745_n400# a_545_n464# a_487_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X18 a_2035_n400# a_1835_n464# a_1777_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X19 a_4099_n400# a_3899_n464# a_3841_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X20 a_n2609_n400# a_n2809_n464# a_n2867_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X21 a_1777_n400# a_1577_n464# a_1519_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X22 a_3841_n400# a_3641_n464# a_3583_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X23 a_n4415_n400# a_n4615_n464# a_n4673_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X24 a_1261_n400# a_1061_n464# a_1003_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X25 a_3583_n400# a_3383_n464# a_3325_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X26 a_n4157_n400# a_n4357_n464# a_n4415_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X27 a_n3899_n400# a_n4099_n464# a_n4157_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X28 a_n1835_n400# a_n2035_n464# a_n2093_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X29 a_2809_n400# a_2609_n464# a_2551_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X30 a_n2351_n400# a_n2551_n464# a_n2609_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X31 a_4357_n400# a_4157_n464# a_4099_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X32 a_4615_n400# a_4415_n464# a_4357_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X33 a_n2093_n400# a_n2293_n464# a_n2351_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X34 a_n29_n400# a_n229_n464# a_n287_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X35 a_229_n400# a_29_n464# a_n29_n400# w_n4873_n697# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
C0 a_n4673_n400# a_n4415_n400# 0.219309f
C1 a_1835_n464# w_n4873_n697# 0.307639f
C2 a_n2867_n400# a_n2609_n400# 0.219309f
C3 a_n2867_n400# a_n3125_n400# 0.219309f
C4 a_4357_n400# a_4099_n400# 0.219309f
C5 a_n3325_n464# w_n4873_n697# 0.307639f
C6 a_3383_n464# w_n4873_n697# 0.307639f
C7 a_803_n464# w_n4873_n697# 0.307639f
C8 a_n1261_n464# w_n4873_n697# 0.307639f
C9 a_n287_n400# a_n545_n400# 0.219309f
C10 a_2035_n400# a_1777_n400# 0.219309f
C11 a_487_n400# a_745_n400# 0.219309f
C12 a_n487_n464# w_n4873_n697# 0.307639f
C13 a_n3641_n400# a_n3899_n400# 0.219309f
C14 a_3899_n464# w_n4873_n697# 0.307639f
C15 a_n29_n400# a_n287_n400# 0.219309f
C16 a_3841_n400# a_3583_n400# 0.219309f
C17 a_n1003_n464# w_n4873_n697# 0.307639f
C18 a_1519_n400# a_1777_n400# 0.219309f
C19 a_n3641_n400# a_n3383_n400# 0.219309f
C20 a_2093_n464# w_n4873_n697# 0.307639f
C21 a_n2351_n400# a_n2609_n400# 0.219309f
C22 w_n4873_n697# a_n3841_n464# 0.307639f
C23 a_n1777_n464# w_n4873_n697# 0.307639f
C24 w_n4873_n697# a_n4615_n464# 0.34286f
C25 a_2035_n400# a_2293_n400# 0.219309f
C26 a_545_n464# w_n4873_n697# 0.307639f
C27 a_1577_n464# w_n4873_n697# 0.307639f
C28 a_4615_n400# w_n4873_n697# 0.249341f
C29 a_1519_n400# a_1261_n400# 0.219309f
C30 a_2351_n464# w_n4873_n697# 0.307639f
C31 a_n745_n464# w_n4873_n697# 0.307639f
C32 a_3841_n400# a_4099_n400# 0.219309f
C33 a_n545_n400# a_n803_n400# 0.219309f
C34 a_745_n400# a_1003_n400# 0.219309f
C35 a_n4673_n400# w_n4873_n697# 0.249341f
C36 a_3641_n464# w_n4873_n697# 0.307639f
C37 a_29_n464# w_n4873_n697# 0.307639f
C38 a_n3067_n464# w_n4873_n697# 0.307639f
C39 a_n1577_n400# a_n1835_n400# 0.219309f
C40 a_3325_n400# a_3583_n400# 0.219309f
C41 a_487_n400# a_229_n400# 0.219309f
C42 w_n4873_n697# a_n4099_n464# 0.307639f
C43 a_n803_n400# a_n1061_n400# 0.219309f
C44 a_n2035_n464# w_n4873_n697# 0.307639f
C45 a_n4157_n400# a_n4415_n400# 0.219309f
C46 a_n2293_n464# w_n4873_n697# 0.307639f
C47 a_2609_n464# w_n4873_n697# 0.307639f
C48 a_287_n464# w_n4873_n697# 0.307639f
C49 a_n229_n464# w_n4873_n697# 0.307639f
C50 a_2551_n400# a_2293_n400# 0.219309f
C51 a_n1061_n400# a_n1319_n400# 0.219309f
C52 a_4615_n400# a_4357_n400# 0.219309f
C53 a_n3383_n400# a_n3125_n400# 0.219309f
C54 w_n4873_n697# a_n1519_n464# 0.307639f
C55 a_3067_n400# a_3325_n400# 0.219309f
C56 a_3125_n464# w_n4873_n697# 0.307639f
C57 a_1261_n400# a_1003_n400# 0.219309f
C58 a_4415_n464# w_n4873_n697# 0.34286f
C59 a_1061_n464# w_n4873_n697# 0.307639f
C60 a_3067_n400# a_2809_n400# 0.219309f
C61 a_1319_n464# w_n4873_n697# 0.307639f
C62 a_n2551_n464# w_n4873_n697# 0.307639f
C63 a_n2809_n464# w_n4873_n697# 0.307639f
C64 a_n2093_n400# a_n2351_n400# 0.219309f
C65 a_n29_n400# a_229_n400# 0.219309f
C66 w_n4873_n697# a_n3583_n464# 0.307639f
C67 a_n2093_n400# a_n1835_n400# 0.219309f
C68 a_2867_n464# w_n4873_n697# 0.307639f
C69 a_4157_n464# w_n4873_n697# 0.307639f
C70 a_n1577_n400# a_n1319_n400# 0.219309f
C71 w_n4873_n697# a_n4357_n464# 0.307639f
C72 a_2551_n400# a_2809_n400# 0.219309f
C73 a_n3899_n400# a_n4157_n400# 0.219309f
C74 a_4615_n400# 0 0.201515f
C75 a_4357_n400# 0 0.116864f
C76 a_4099_n400# 0 0.116864f
C77 a_3841_n400# 0 0.116864f
C78 a_3583_n400# 0 0.116864f
C79 a_3325_n400# 0 0.116864f
C80 a_3067_n400# 0 0.116864f
C81 a_2809_n400# 0 0.116864f
C82 a_2551_n400# 0 0.116864f
C83 a_2293_n400# 0 0.116864f
C84 a_2035_n400# 0 0.116864f
C85 a_1777_n400# 0 0.116864f
C86 a_1519_n400# 0 0.116864f
C87 a_1261_n400# 0 0.116864f
C88 a_1003_n400# 0 0.116864f
C89 a_745_n400# 0 0.116864f
C90 a_487_n400# 0 0.116864f
C91 a_229_n400# 0 0.116864f
C92 a_n29_n400# 0 0.116864f
C93 a_n287_n400# 0 0.116864f
C94 a_n545_n400# 0 0.116864f
C95 a_n803_n400# 0 0.116864f
C96 a_n1061_n400# 0 0.116864f
C97 a_n1319_n400# 0 0.116864f
C98 a_n1577_n400# 0 0.116864f
C99 a_n1835_n400# 0 0.116864f
C100 a_n2093_n400# 0 0.116864f
C101 a_n2351_n400# 0 0.116864f
C102 a_n2609_n400# 0 0.116864f
C103 a_n2867_n400# 0 0.116864f
C104 a_n3125_n400# 0 0.116864f
C105 a_n3383_n400# 0 0.116864f
C106 a_n3641_n400# 0 0.116864f
C107 a_n3899_n400# 0 0.116864f
C108 a_n4157_n400# 0 0.116864f
C109 a_n4415_n400# 0 0.116864f
C110 a_n4673_n400# 0 0.201515f
C111 a_4415_n464# 0 0.233871f
C112 a_4157_n464# 0 0.211442f
C113 a_3899_n464# 0 0.211442f
C114 a_3641_n464# 0 0.211442f
C115 a_3383_n464# 0 0.211442f
C116 a_3125_n464# 0 0.211442f
C117 a_2867_n464# 0 0.211442f
C118 a_2609_n464# 0 0.211442f
C119 a_2351_n464# 0 0.211442f
C120 a_2093_n464# 0 0.211442f
C121 a_1835_n464# 0 0.211442f
C122 a_1577_n464# 0 0.211442f
C123 a_1319_n464# 0 0.211442f
C124 a_1061_n464# 0 0.211442f
C125 a_803_n464# 0 0.211442f
C126 a_545_n464# 0 0.211442f
C127 a_287_n464# 0 0.211442f
C128 a_29_n464# 0 0.211442f
C129 a_n229_n464# 0 0.211442f
C130 a_n487_n464# 0 0.211442f
C131 a_n745_n464# 0 0.211442f
C132 a_n1003_n464# 0 0.211442f
C133 a_n1261_n464# 0 0.211442f
C134 a_n1519_n464# 0 0.211442f
C135 a_n1777_n464# 0 0.211442f
C136 a_n2035_n464# 0 0.211442f
C137 a_n2293_n464# 0 0.211442f
C138 a_n2551_n464# 0 0.211442f
C139 a_n2809_n464# 0 0.211442f
C140 a_n3067_n464# 0 0.211442f
C141 a_n3325_n464# 0 0.211442f
C142 a_n3583_n464# 0 0.211442f
C143 a_n3841_n464# 0 0.211442f
C144 a_n4099_n464# 0 0.211442f
C145 a_n4357_n464# 0 0.211442f
C146 a_n4615_n464# 0 0.233871f
C147 w_n4873_n697# 0 47.096104f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_Z5XS7R c1_6184_n8000# c1_n8876_n8000# m3_6144_n8040#
+ c1_160_n8000# m3_n2892_n8040# m3_n8916_n8040# c1_3172_n8000# c1_n5864_n8000# m3_3132_n8040#
+ m3_n5904_n8040# m3_120_n8040# c1_n2852_n8000#
X0 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X1 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X2 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X3 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X4 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X5 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X6 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X7 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X8 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X9 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X10 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X11 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X12 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X13 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X14 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X15 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X16 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X17 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X18 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X19 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X20 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X21 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X22 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X23 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X24 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X25 c1_n8876_n8000# m3_n8916_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X26 c1_6184_n8000# m3_6144_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X27 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X28 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X29 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X30 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X31 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 c1_160_n8000# m3_120_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X33 c1_3172_n8000# m3_3132_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 c1_n5864_n8000# m3_n5904_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X35 c1_n2852_n8000# m3_n2892_n8040# sky130_fd_pr__cap_mim_m3_1 l=12 w=12
C0 m3_n2892_n8040# c1_160_n8000# 3.17007f
C1 m3_3132_n8040# m3_120_n8040# 3.84418f
C2 m3_n2892_n8040# m3_n5904_n8040# 3.84418f
C3 c1_n2852_n8000# m3_n2892_n8040# 81.8286f
C4 c1_3172_n8000# m3_3132_n8040# 81.8286f
C5 m3_6144_n8040# c1_6184_n8000# 81.8286f
C6 c1_n2852_n8000# m3_n5904_n8040# 3.17007f
C7 c1_160_n8000# m3_120_n8040# 81.8286f
C8 m3_n2892_n8040# m3_120_n8040# 3.84418f
C9 c1_n5864_n8000# m3_n5904_n8040# 81.8286f
C10 m3_n8916_n8040# m3_n5904_n8040# 3.84418f
C11 m3_6144_n8040# m3_3132_n8040# 3.84418f
C12 c1_3172_n8000# m3_120_n8040# 3.17007f
C13 m3_n8916_n8040# c1_n5864_n8000# 3.17007f
C14 m3_n8916_n8040# c1_n8876_n8000# 81.8286f
C15 c1_6184_n8000# m3_3132_n8040# 3.17007f
C16 c1_6184_n8000# 0 1.97709f
C17 c1_3172_n8000# 0 1.97709f
C18 c1_160_n8000# 0 1.97709f
C19 c1_n2852_n8000# 0 1.97709f
C20 c1_n5864_n8000# 0 1.97709f
C21 c1_n8876_n8000# 0 4.298831f
C22 m3_6144_n8040# 0 21.7528f
C23 m3_3132_n8040# 0 16.7642f
C24 m3_120_n8040# 0 16.7642f
C25 m3_n2892_n8040# 0 16.7642f
C26 m3_n5904_n8040# 0 16.7642f
C27 m3_n8916_n8040# 0 19.2536f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_EVM3FM a_29_n964# a_n129_n964# a_187_n964# a_445_n900#
+ a_n287_n964# a_345_n964# a_603_n900# a_n445_n964# a_761_n900# a_503_n964# a_n29_n900#
+ a_n603_n964# a_661_n964# a_n187_n900# a_n761_n964# a_n819_n900# a_n345_n900# a_129_n900#
+ a_n503_n900# w_n1019_n1197# a_n661_n900# a_287_n900#
X0 a_n187_n900# a_n287_n964# a_n345_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X1 a_761_n900# a_661_n964# a_603_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=0.5
X2 a_287_n900# a_187_n964# a_129_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X3 a_n345_n900# a_n445_n964# a_n503_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X4 a_129_n900# a_29_n964# a_n29_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X5 a_445_n900# a_345_n964# a_287_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X6 a_n503_n900# a_n603_n964# a_n661_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X7 a_n29_n900# a_n129_n964# a_n187_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X8 a_603_n900# a_503_n964# a_445_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=0.5
X9 a_n661_n900# a_n761_n964# a_n819_n900# w_n1019_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=0.5
C0 w_n1019_n1197# a_187_n964# 0.180946f
C1 a_603_n900# a_661_n964# 0.115387f
C2 a_n503_n900# a_n445_n964# 0.115387f
C3 a_n761_n964# a_n819_n900# 0.115387f
C4 a_445_n900# a_603_n900# 0.801423f
C5 a_n29_n900# a_n129_n964# 0.115387f
C6 a_445_n900# a_287_n900# 0.801423f
C7 a_129_n900# a_187_n964# 0.115387f
C8 a_n503_n900# a_n661_n900# 0.801423f
C9 w_n1019_n1197# a_n761_n964# 0.220136f
C10 a_n29_n900# a_n187_n900# 0.801423f
C11 a_n345_n900# a_n287_n964# 0.115387f
C12 a_n29_n900# a_129_n900# 0.801423f
C13 a_345_n964# a_287_n900# 0.115387f
C14 w_n1019_n1197# a_n819_n900# 0.529882f
C15 a_761_n900# a_603_n900# 0.801423f
C16 a_n503_n900# a_n603_n964# 0.115387f
C17 w_n1019_n1197# a_n129_n964# 0.180946f
C18 w_n1019_n1197# a_n287_n964# 0.180946f
C19 a_n345_n900# a_n187_n900# 0.801423f
C20 a_n187_n900# a_n129_n964# 0.115387f
C21 a_n287_n964# a_n187_n900# 0.115387f
C22 a_287_n900# a_187_n964# 0.115387f
C23 a_761_n900# a_661_n964# 0.115387f
C24 a_n345_n900# a_n445_n964# 0.115387f
C25 a_n761_n964# a_n661_n900# 0.115387f
C26 a_345_n964# a_445_n900# 0.115387f
C27 w_n1019_n1197# a_503_n964# 0.180946f
C28 a_29_n964# a_n29_n900# 0.115387f
C29 w_n1019_n1197# a_n445_n964# 0.180946f
C30 a_n661_n900# a_n819_n900# 0.801423f
C31 a_29_n964# w_n1019_n1197# 0.180946f
C32 a_603_n900# a_503_n964# 0.115387f
C33 w_n1019_n1197# a_n603_n964# 0.180946f
C34 a_29_n964# a_129_n900# 0.115387f
C35 w_n1019_n1197# a_661_n964# 0.220136f
C36 a_129_n900# a_287_n900# 0.801423f
C37 a_445_n900# a_503_n964# 0.115387f
C38 a_n345_n900# a_n503_n900# 0.801423f
C39 a_n603_n964# a_n661_n900# 0.115387f
C40 w_n1019_n1197# a_345_n964# 0.180946f
C41 w_n1019_n1197# a_761_n900# 0.529882f
C42 a_761_n900# 0 0.393686f
C43 a_603_n900# 0 0.155127f
C44 a_445_n900# 0 0.155127f
C45 a_287_n900# 0 0.155127f
C46 a_129_n900# 0 0.155127f
C47 a_n29_n900# 0 0.155127f
C48 a_n187_n900# 0 0.155127f
C49 a_n345_n900# 0 0.155127f
C50 a_n503_n900# 0 0.155127f
C51 a_n661_n900# 0 0.155127f
C52 a_n819_n900# 0 0.393686f
C53 a_661_n964# 0 0.135226f
C54 a_503_n964# 0 0.112152f
C55 a_345_n964# 0 0.112152f
C56 a_187_n964# 0 0.112152f
C57 a_29_n964# 0 0.112152f
C58 a_n129_n964# 0 0.112152f
C59 a_n287_n964# 0 0.112152f
C60 a_n445_n964# 0 0.112152f
C61 a_n603_n964# 0 0.112152f
C62 a_n761_n964# 0 0.135226f
C63 w_n1019_n1197# 0 16.885199f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN a_n2093_n200# a_803_n255# a_n2035_n255#
+ a_n3841_n255# a_1261_n200# a_n4357_n255# a_3583_n200# a_n1319_n200# a_n4415_n200#
+ a_3125_n255# a_1835_n255# a_n287_n200# a_n229_n255# a_4099_n200# a_n1061_n200# a_287_n255#
+ a_n1003_n255# a_2809_n200# a_745_n200# a_n3383_n200# a_2093_n255# a_n3325_n255#
+ a_2551_n200# a_3067_n200# a_4415_n255# a_1319_n255# a_4873_n200# a_1777_n200# a_n2609_n200#
+ a_n2293_n255# a_1061_n255# a_n2351_n200# a_229_n200# a_3383_n255# a_n1577_n200#
+ a_n4673_n200# a_n1519_n255# a_n4615_n255# a_3841_n200# a_2035_n200# a_n487_n255#
+ a_n545_n200# a_n3899_n200# a_n1261_n255# a_4357_n200# a_2609_n255# a_545_n255# a_n3583_n255#
+ a_n3641_n200# a_2351_n255# a_1003_n200# a_n4099_n255# a_n4157_n200# a_4673_n255#
+ a_1577_n255# a_3325_n200# a_n2867_n200# a_n2809_n255# a_3899_n255# a_n2551_n255#
+ a_487_n200# a_n29_n200# a_n3067_n255# a_2293_n200# a_29_n255# a_n1777_n255# a_n4873_n255#
+ a_n1835_n200# a_n3125_n200# a_n4931_n200# a_3641_n255# a_4157_n255# a_n745_n255#
+ a_n803_n200# a_2867_n255# a_4615_n200# a_1519_n200# a_n5065_n422#
X0 a_487_n200# a_287_n255# a_229_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_2035_n200# a_1835_n255# a_1777_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_4099_n200# a_3899_n255# a_3841_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_n2609_n200# a_n2809_n255# a_n2867_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_1777_n200# a_1577_n255# a_1519_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_3841_n200# a_3641_n255# a_3583_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n4415_n200# a_n4615_n255# a_n4673_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_1261_n200# a_1061_n255# a_1003_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_3583_n200# a_3383_n255# a_3325_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n4157_n200# a_n4357_n255# a_n4415_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n3899_n200# a_n4099_n255# a_n4157_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1835_n200# a_n2035_n255# a_n2093_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X12 a_n4673_n200# a_n4873_n255# a_n4931_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X13 a_2809_n200# a_2609_n255# a_2551_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X14 a_n2351_n200# a_n2551_n255# a_n2609_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X15 a_4357_n200# a_4157_n255# a_4099_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X16 a_4615_n200# a_4415_n255# a_4357_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X17 a_n2093_n200# a_n2293_n255# a_n2351_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X18 a_n29_n200# a_n229_n255# a_n287_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X19 a_229_n200# a_29_n255# a_n29_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X20 a_3067_n200# a_2867_n255# a_2809_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X21 a_4873_n200# a_4673_n255# a_4615_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X22 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X23 a_n545_n200# a_n745_n255# a_n803_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X24 a_2293_n200# a_2093_n255# a_2035_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X25 a_2551_n200# a_2351_n255# a_2293_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X26 a_n3125_n200# a_n3325_n255# a_n3383_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X27 a_n2867_n200# a_n3067_n255# a_n3125_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X28 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X29 a_n287_n200# a_n487_n255# a_n545_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X30 a_n3641_n200# a_n3841_n255# a_n3899_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X31 a_n1577_n200# a_n1777_n255# a_n1835_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X32 a_1519_n200# a_1319_n255# a_1261_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X33 a_n3383_n200# a_n3583_n255# a_n3641_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X34 a_3325_n200# a_3125_n255# a_3067_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X35 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X36 a_745_n200# a_545_n255# a_487_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X37 a_1003_n200# a_803_n255# a_745_n200# a_n5065_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
C0 a_3325_n200# a_3583_n200# 0.110175f
C1 a_n2609_n200# a_n2867_n200# 0.110175f
C2 a_n3125_n200# a_n2867_n200# 0.110175f
C3 a_2293_n200# a_2551_n200# 0.110175f
C4 a_n1061_n200# a_n1319_n200# 0.110175f
C5 a_1261_n200# a_1003_n200# 0.110175f
C6 a_n4157_n200# a_n3899_n200# 0.110175f
C7 a_n287_n200# a_n29_n200# 0.110175f
C8 a_3325_n200# a_3067_n200# 0.110175f
C9 a_n3125_n200# a_n3383_n200# 0.110175f
C10 a_1261_n200# a_1519_n200# 0.110175f
C11 a_3841_n200# a_3583_n200# 0.110175f
C12 a_n1061_n200# a_n803_n200# 0.110175f
C13 a_4099_n200# a_3841_n200# 0.110175f
C14 a_n545_n200# a_n803_n200# 0.110175f
C15 a_2551_n200# a_2809_n200# 0.110175f
C16 a_n287_n200# a_n545_n200# 0.110175f
C17 a_n4415_n200# a_n4157_n200# 0.110175f
C18 a_4615_n200# a_4357_n200# 0.110175f
C19 a_n3641_n200# a_n3383_n200# 0.110175f
C20 a_229_n200# a_n29_n200# 0.110175f
C21 a_n1577_n200# a_n1319_n200# 0.110175f
C22 a_2293_n200# a_2035_n200# 0.110175f
C23 a_1003_n200# a_745_n200# 0.110175f
C24 a_4099_n200# a_4357_n200# 0.110175f
C25 a_n3899_n200# a_n3641_n200# 0.110175f
C26 a_n2351_n200# a_n2093_n200# 0.110175f
C27 a_1777_n200# a_1519_n200# 0.110175f
C28 a_745_n200# a_487_n200# 0.110175f
C29 a_n4415_n200# a_n4673_n200# 0.110175f
C30 a_n1835_n200# a_n1577_n200# 0.110175f
C31 a_3067_n200# a_2809_n200# 0.110175f
C32 a_n2351_n200# a_n2609_n200# 0.110175f
C33 a_n1835_n200# a_n2093_n200# 0.110175f
C34 a_1777_n200# a_2035_n200# 0.110175f
C35 a_n4931_n200# a_n4673_n200# 0.110175f
C36 a_4873_n200# a_4615_n200# 0.110175f
C37 a_229_n200# a_487_n200# 0.110175f
C38 a_4873_n200# a_n5065_n422# 0.241444f
C39 a_n4931_n200# a_n5065_n422# 0.241444f
C40 a_4673_n255# a_n5065_n422# 0.55256f
C41 a_4415_n255# a_n5065_n422# 0.498389f
C42 a_4157_n255# a_n5065_n422# 0.498389f
C43 a_3899_n255# a_n5065_n422# 0.498389f
C44 a_3641_n255# a_n5065_n422# 0.498389f
C45 a_3383_n255# a_n5065_n422# 0.498389f
C46 a_3125_n255# a_n5065_n422# 0.498389f
C47 a_2867_n255# a_n5065_n422# 0.498389f
C48 a_2609_n255# a_n5065_n422# 0.498389f
C49 a_2351_n255# a_n5065_n422# 0.498389f
C50 a_2093_n255# a_n5065_n422# 0.498389f
C51 a_1835_n255# a_n5065_n422# 0.498389f
C52 a_1577_n255# a_n5065_n422# 0.498389f
C53 a_1319_n255# a_n5065_n422# 0.498389f
C54 a_1061_n255# a_n5065_n422# 0.498389f
C55 a_803_n255# a_n5065_n422# 0.498389f
C56 a_545_n255# a_n5065_n422# 0.498389f
C57 a_287_n255# a_n5065_n422# 0.498389f
C58 a_29_n255# a_n5065_n422# 0.498389f
C59 a_n229_n255# a_n5065_n422# 0.498389f
C60 a_n487_n255# a_n5065_n422# 0.498389f
C61 a_n745_n255# a_n5065_n422# 0.498389f
C62 a_n1003_n255# a_n5065_n422# 0.498389f
C63 a_n1261_n255# a_n5065_n422# 0.498389f
C64 a_n1519_n255# a_n5065_n422# 0.498389f
C65 a_n1777_n255# a_n5065_n422# 0.498389f
C66 a_n2035_n255# a_n5065_n422# 0.498389f
C67 a_n2293_n255# a_n5065_n422# 0.498389f
C68 a_n2551_n255# a_n5065_n422# 0.498389f
C69 a_n2809_n255# a_n5065_n422# 0.498389f
C70 a_n3067_n255# a_n5065_n422# 0.498389f
C71 a_n3325_n255# a_n5065_n422# 0.498389f
C72 a_n3583_n255# a_n5065_n422# 0.498389f
C73 a_n3841_n255# a_n5065_n422# 0.498389f
C74 a_n4099_n255# a_n5065_n422# 0.498389f
C75 a_n4357_n255# a_n5065_n422# 0.498389f
C76 a_n4615_n255# a_n5065_n422# 0.498389f
C77 a_n4873_n255# a_n5065_n422# 0.55256f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_Q46EE6 a_1261_n200# a_n487_n264# a_n1261_n264#
+ w_n2035_n497# a_n1319_n200# a_545_n264# a_n287_n200# a_n1061_n200# a_1577_n264#
+ a_745_n200# a_1777_n200# a_n1777_n264# a_29_n264# a_229_n200# a_n745_n264# a_n1577_n200#
+ a_803_n264# a_n545_n200# a_1003_n200# a_n229_n264# a_n1003_n264# a_287_n264# a_487_n200#
+ a_n29_n200# a_1319_n264# a_n1835_n200# a_1061_n264# a_n803_n200# a_1519_n200# a_n1519_n264#
X0 a_745_n200# a_545_n264# a_487_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1003_n200# a_803_n264# a_745_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_487_n200# a_287_n264# a_229_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_1777_n200# a_1577_n264# a_1519_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X4 a_1261_n200# a_1061_n264# a_1003_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X5 a_n29_n200# a_n229_n264# a_n287_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_229_n200# a_29_n264# a_n29_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n1319_n200# a_n1519_n264# a_n1577_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_n545_n200# a_n745_n264# a_n803_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X9 a_n803_n200# a_n1003_n264# a_n1061_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_n287_n200# a_n487_n264# a_n545_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_n1577_n200# a_n1777_n264# a_n1835_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X12 a_1519_n200# a_1319_n264# a_1261_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X13 a_n1061_n200# a_n1261_n264# a_n1319_n200# w_n2035_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
C0 a_1061_n264# w_n2035_n497# 0.307639f
C1 a_n745_n264# w_n2035_n497# 0.307639f
C2 a_n29_n200# a_229_n200# 0.110175f
C3 a_n1519_n264# w_n2035_n497# 0.307639f
C4 a_29_n264# w_n2035_n497# 0.307639f
C5 a_1003_n200# a_745_n200# 0.110175f
C6 a_287_n264# w_n2035_n497# 0.307639f
C7 a_487_n200# a_745_n200# 0.110175f
C8 a_n1835_n200# w_n2035_n497# 0.137129f
C9 a_803_n264# w_n2035_n497# 0.307639f
C10 a_n1577_n200# a_n1835_n200# 0.110175f
C11 a_1577_n264# w_n2035_n497# 0.34286f
C12 a_n29_n200# a_n287_n200# 0.110175f
C13 a_n803_n200# a_n545_n200# 0.110175f
C14 a_n487_n264# w_n2035_n497# 0.307639f
C15 a_1777_n200# w_n2035_n497# 0.137129f
C16 a_487_n200# a_229_n200# 0.110175f
C17 a_n1777_n264# w_n2035_n497# 0.34286f
C18 a_n1577_n200# a_n1319_n200# 0.110175f
C19 a_545_n264# w_n2035_n497# 0.307639f
C20 a_n1061_n200# a_n1319_n200# 0.110175f
C21 a_n803_n200# a_n1061_n200# 0.110175f
C22 a_1319_n264# w_n2035_n497# 0.307639f
C23 a_n229_n264# w_n2035_n497# 0.307639f
C24 a_n287_n200# a_n545_n200# 0.110175f
C25 a_n1261_n264# w_n2035_n497# 0.307639f
C26 a_1261_n200# a_1519_n200# 0.110175f
C27 a_1261_n200# a_1003_n200# 0.110175f
C28 a_1777_n200# a_1519_n200# 0.110175f
C29 a_n1003_n264# w_n2035_n497# 0.307639f
C30 a_1777_n200# 0 0.104989f
C31 a_n1835_n200# 0 0.104989f
C32 a_1577_n264# 0 0.227252f
C33 a_1319_n264# 0 0.204823f
C34 a_1061_n264# 0 0.204823f
C35 a_803_n264# 0 0.204823f
C36 a_545_n264# 0 0.204823f
C37 a_287_n264# 0 0.204823f
C38 a_29_n264# 0 0.204823f
C39 a_n229_n264# 0 0.204823f
C40 a_n487_n264# 0 0.204823f
C41 a_n745_n264# 0 0.204823f
C42 a_n1003_n264# 0 0.204823f
C43 a_n1261_n264# 0 0.204823f
C44 a_n1519_n264# 0 0.204823f
C45 a_n1777_n264# 0 0.227252f
C46 w_n2035_n497# 0 14.831599f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_UGZTXE a_1061_n655# a_n2293_n655# a_n2351_n600#
+ a_229_n600# a_n1577_n600# a_3383_n655# a_n1519_n655# a_2035_n600# a_n487_n655# a_n1261_n655#
+ a_n545_n600# a_2609_n655# a_545_n655# a_2351_n655# a_n3583_n655# a_1003_n600# a_n3641_n600#
+ a_1577_n655# a_n2867_n600# a_n2809_n655# a_3325_n600# a_n2551_n655# a_n29_n600#
+ a_487_n600# a_n1777_n655# a_n3067_n655# a_2293_n600# a_n3125_n600# a_29_n655# a_n1835_n600#
+ a_2867_n655# a_n745_n655# a_n803_n600# a_1519_n600# a_n2093_n600# a_803_n655# a_n2035_n655#
+ a_n3775_n822# a_1261_n600# a_3125_n655# a_3583_n600# a_n1319_n600# a_1835_n655#
+ a_n287_n600# a_n1061_n600# a_n229_n655# a_n1003_n655# a_287_n655# a_2809_n600# a_2093_n655#
+ a_745_n600# a_n3383_n600# a_n3325_n655# a_2551_n600# a_3067_n600# a_1777_n600# a_n2609_n600#
+ a_1319_n655#
X0 a_2809_n600# a_2609_n655# a_2551_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X1 a_n2351_n600# a_n2551_n655# a_n2609_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X2 a_n2093_n600# a_n2293_n655# a_n2351_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X3 a_229_n600# a_29_n655# a_n29_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X4 a_n29_n600# a_n229_n655# a_n287_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X5 a_3067_n600# a_2867_n655# a_2809_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X6 a_n1319_n600# a_n1519_n655# a_n1577_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X7 a_2551_n600# a_2351_n655# a_2293_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X8 a_n3125_n600# a_n3325_n655# a_n3383_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X9 a_n545_n600# a_n745_n655# a_n803_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X10 a_n287_n600# a_n487_n655# a_n545_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X11 a_2293_n600# a_2093_n655# a_2035_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X12 a_n2867_n600# a_n3067_n655# a_n3125_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X13 a_n803_n600# a_n1003_n655# a_n1061_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X14 a_n3383_n600# a_n3583_n655# a_n3641_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.58 w=6 l=1
X15 a_n1577_n600# a_n1777_n655# a_n1835_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X16 a_1519_n600# a_1319_n655# a_1261_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X17 a_n1061_n600# a_n1261_n655# a_n1319_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X18 a_3325_n600# a_3125_n655# a_3067_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X19 a_1003_n600# a_803_n655# a_745_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X20 a_745_n600# a_545_n655# a_487_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X21 a_487_n600# a_287_n655# a_229_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X22 a_2035_n600# a_1835_n655# a_1777_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X23 a_n2609_n600# a_n2809_n655# a_n2867_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X24 a_1777_n600# a_1577_n655# a_1519_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X25 a_3583_n600# a_3383_n655# a_3325_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.58 as=0.87 ps=6.29 w=6 l=1
X26 a_1261_n600# a_1061_n655# a_1003_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
X27 a_n1835_n600# a_n2035_n655# a_n2093_n600# a_n3775_n822# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=1
C0 a_n2867_n600# a_n2609_n600# 0.328443f
C1 a_n2351_n600# a_n2551_n655# 0.133664f
C2 a_487_n600# a_229_n600# 0.328443f
C3 a_3125_n655# a_3325_n600# 0.133664f
C4 a_2609_n655# a_2809_n600# 0.133664f
C5 a_1519_n600# a_1577_n655# 0.133664f
C6 a_n1577_n600# a_n1777_n655# 0.133664f
C7 a_n1319_n600# a_n1261_n655# 0.133664f
C8 a_1061_n655# a_1003_n600# 0.133664f
C9 a_n3641_n600# a_n3583_n655# 0.133664f
C10 a_29_n655# a_229_n600# 0.133664f
C11 a_2293_n600# a_2035_n600# 0.328443f
C12 a_n1061_n600# a_n1003_n655# 0.133664f
C13 a_n803_n600# a_n1003_n655# 0.133664f
C14 a_287_n655# a_229_n600# 0.133664f
C15 a_1003_n600# a_745_n600# 0.328443f
C16 a_n2867_n600# a_n3125_n600# 0.328443f
C17 a_2293_n600# a_2551_n600# 0.328443f
C18 a_1777_n600# a_1519_n600# 0.328443f
C19 a_n3383_n600# a_n3125_n600# 0.328443f
C20 a_n2809_n655# a_n2867_n600# 0.133664f
C21 a_n2351_n600# a_n2609_n600# 0.328443f
C22 a_n545_n600# a_n803_n600# 0.328443f
C23 a_1519_n600# a_1319_n655# 0.133664f
C24 a_2293_n600# a_2351_n655# 0.133664f
C25 a_n287_n600# a_n487_n655# 0.133664f
C26 a_n545_n600# a_n487_n655# 0.133664f
C27 a_2293_n600# a_2093_n655# 0.133664f
C28 a_3383_n655# a_3583_n600# 0.133664f
C29 a_1319_n655# a_1261_n600# 0.133664f
C30 a_n1061_n600# a_n1319_n600# 0.328443f
C31 a_1061_n655# a_1261_n600# 0.133664f
C32 a_545_n655# a_745_n600# 0.133664f
C33 a_n1835_n600# a_n1777_n655# 0.133664f
C34 a_3067_n600# a_3325_n600# 0.328443f
C35 a_n3125_n600# a_n3325_n655# 0.133664f
C36 a_1003_n600# a_1261_n600# 0.328443f
C37 a_487_n600# a_745_n600# 0.328443f
C38 a_n2551_n655# a_n2609_n600# 0.133664f
C39 a_n29_n600# a_n229_n655# 0.133664f
C40 a_1003_n600# a_803_n655# 0.133664f
C41 a_803_n655# a_745_n600# 0.133664f
C42 a_n2093_n600# a_n2035_n655# 0.133664f
C43 a_n287_n600# a_n229_n655# 0.133664f
C44 a_n1577_n600# a_n1519_n655# 0.133664f
C45 a_n2093_n600# a_n1835_n600# 0.328443f
C46 a_n745_n655# a_n803_n600# 0.133664f
C47 a_2035_n600# a_1835_n655# 0.133664f
C48 a_3325_n600# a_3583_n600# 0.328443f
C49 a_3067_n600# a_3125_n655# 0.133664f
C50 a_n29_n600# a_n287_n600# 0.328443f
C51 a_n3383_n600# a_n3325_n655# 0.133664f
C52 a_2035_n600# a_2093_n655# 0.133664f
C53 a_n3641_n600# a_n3383_n600# 0.328443f
C54 a_n545_n600# a_n287_n600# 0.328443f
C55 a_2551_n600# a_2351_n655# 0.133664f
C56 a_1519_n600# a_1261_n600# 0.328443f
C57 a_n1319_n600# a_n1577_n600# 0.328443f
C58 a_545_n655# a_487_n600# 0.133664f
C59 a_n1061_n600# a_n1261_n655# 0.133664f
C60 a_1777_n600# a_2035_n600# 0.328443f
C61 a_n2293_n655# a_n2351_n600# 0.133664f
C62 a_n1319_n600# a_n1519_n655# 0.133664f
C63 a_n1577_n600# a_n1835_n600# 0.328443f
C64 a_29_n655# a_n29_n600# 0.133664f
C65 a_2551_n600# a_2809_n600# 0.328443f
C66 a_n2293_n655# a_n2093_n600# 0.133664f
C67 a_1777_n600# a_1835_n655# 0.133664f
C68 a_1777_n600# a_1577_n655# 0.133664f
C69 a_3383_n655# a_3325_n600# 0.133664f
C70 a_n3067_n655# a_n3125_n600# 0.133664f
C71 a_n545_n600# a_n745_n655# 0.133664f
C72 a_287_n655# a_487_n600# 0.133664f
C73 a_2551_n600# a_2609_n655# 0.133664f
C74 a_3067_n600# a_2867_n655# 0.133664f
C75 a_n2351_n600# a_n2093_n600# 0.328443f
C76 a_3067_n600# a_2809_n600# 0.328443f
C77 a_n3067_n655# a_n2867_n600# 0.133664f
C78 a_n2809_n655# a_n2609_n600# 0.133664f
C79 a_n1061_n600# a_n803_n600# 0.328443f
C80 a_2867_n655# a_2809_n600# 0.133664f
C81 a_n29_n600# a_229_n600# 0.328443f
C82 a_n3583_n655# a_n3383_n600# 0.133664f
C83 a_n1835_n600# a_n2035_n655# 0.133664f
C84 a_3583_n600# a_n3775_n822# 0.657435f
C85 a_3325_n600# a_n3775_n822# 0.193606f
C86 a_3067_n600# a_n3775_n822# 0.193606f
C87 a_2809_n600# a_n3775_n822# 0.193606f
C88 a_2551_n600# a_n3775_n822# 0.193606f
C89 a_2293_n600# a_n3775_n822# 0.193606f
C90 a_2035_n600# a_n3775_n822# 0.193606f
C91 a_1777_n600# a_n3775_n822# 0.193606f
C92 a_1519_n600# a_n3775_n822# 0.193606f
C93 a_1261_n600# a_n3775_n822# 0.193606f
C94 a_1003_n600# a_n3775_n822# 0.193606f
C95 a_745_n600# a_n3775_n822# 0.193606f
C96 a_487_n600# a_n3775_n822# 0.193606f
C97 a_229_n600# a_n3775_n822# 0.193606f
C98 a_n29_n600# a_n3775_n822# 0.193606f
C99 a_n287_n600# a_n3775_n822# 0.193606f
C100 a_n545_n600# a_n3775_n822# 0.193606f
C101 a_n803_n600# a_n3775_n822# 0.193606f
C102 a_n1061_n600# a_n3775_n822# 0.193606f
C103 a_n1319_n600# a_n3775_n822# 0.193606f
C104 a_n1577_n600# a_n3775_n822# 0.193606f
C105 a_n1835_n600# a_n3775_n822# 0.193606f
C106 a_n2093_n600# a_n3775_n822# 0.193606f
C107 a_n2351_n600# a_n3775_n822# 0.193606f
C108 a_n2609_n600# a_n3775_n822# 0.193606f
C109 a_n2867_n600# a_n3775_n822# 0.193606f
C110 a_n3125_n600# a_n3775_n822# 0.193606f
C111 a_n3383_n600# a_n3775_n822# 0.193606f
C112 a_n3641_n600# a_n3775_n822# 0.657435f
C113 a_3383_n655# a_n3775_n822# 0.562598f
C114 a_3125_n655# a_n3775_n822# 0.508426f
C115 a_2867_n655# a_n3775_n822# 0.508426f
C116 a_2609_n655# a_n3775_n822# 0.508426f
C117 a_2351_n655# a_n3775_n822# 0.508426f
C118 a_2093_n655# a_n3775_n822# 0.508426f
C119 a_1835_n655# a_n3775_n822# 0.508426f
C120 a_1577_n655# a_n3775_n822# 0.508426f
C121 a_1319_n655# a_n3775_n822# 0.508426f
C122 a_1061_n655# a_n3775_n822# 0.508426f
C123 a_803_n655# a_n3775_n822# 0.508426f
C124 a_545_n655# a_n3775_n822# 0.508426f
C125 a_287_n655# a_n3775_n822# 0.508426f
C126 a_29_n655# a_n3775_n822# 0.508426f
C127 a_n229_n655# a_n3775_n822# 0.508426f
C128 a_n487_n655# a_n3775_n822# 0.508426f
C129 a_n745_n655# a_n3775_n822# 0.508426f
C130 a_n1003_n655# a_n3775_n822# 0.508426f
C131 a_n1261_n655# a_n3775_n822# 0.508426f
C132 a_n1519_n655# a_n3775_n822# 0.508426f
C133 a_n1777_n655# a_n3775_n822# 0.508426f
C134 a_n2035_n655# a_n3775_n822# 0.508426f
C135 a_n2293_n655# a_n3775_n822# 0.508426f
C136 a_n2551_n655# a_n3775_n822# 0.508426f
C137 a_n2809_n655# a_n3775_n822# 0.508426f
C138 a_n3067_n655# a_n3775_n822# 0.508426f
C139 a_n3325_n655# a_n3775_n822# 0.508426f
C140 a_n3583_n655# a_n3775_n822# 0.562598f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_XW23Q2 a_29_n964# a_n2351_n900# a_229_n900# a_n745_n964#
+ a_n1577_n900# a_2035_n900# a_803_n964# a_n2035_n964# a_n545_n900# a_1835_n964# a_1003_n900#
+ a_n229_n964# a_n1003_n964# a_287_n964# a_n2867_n900# a_2093_n964# a_487_n900# a_n29_n900#
+ a_2293_n900# a_1319_n964# a_n1835_n900# a_1061_n964# a_n2293_n964# a_n803_n900#
+ a_1519_n900# a_n2093_n900# a_n1519_n964# a_1261_n900# a_n487_n964# a_n1261_n964#
+ a_2609_n964# a_n1319_n900# a_545_n964# a_n287_n900# a_2351_n964# a_n1061_n900# a_1577_n964#
+ a_2809_n900# a_745_n900# a_n2809_n964# a_2551_n900# a_n2551_n964# w_n3067_n1197#
+ a_1777_n900# a_n2609_n900# a_n1777_n964#
X0 a_n2609_n900# a_n2809_n964# a_n2867_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=2.61 ps=18.58 w=9 l=1
X1 a_1261_n900# a_1061_n964# a_1003_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X2 a_n1835_n900# a_n2035_n964# a_n2093_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X3 a_2809_n900# a_2609_n964# a_2551_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.61 pd=18.58 as=1.305 ps=9.29 w=9 l=1
X4 a_n2351_n900# a_n2551_n964# a_n2609_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X5 a_n2093_n900# a_n2293_n964# a_n2351_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X6 a_n29_n900# a_n229_n964# a_n287_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X7 a_229_n900# a_29_n964# a_n29_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X8 a_n1319_n900# a_n1519_n964# a_n1577_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X9 a_2551_n900# a_2351_n964# a_2293_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X10 a_n545_n900# a_n745_n964# a_n803_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X11 a_n287_n900# a_n487_n964# a_n545_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X12 a_2293_n900# a_2093_n964# a_2035_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X13 a_n803_n900# a_n1003_n964# a_n1061_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X14 a_n1577_n900# a_n1777_n964# a_n1835_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X15 a_1519_n900# a_1319_n964# a_1261_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X16 a_n1061_n900# a_n1261_n964# a_n1319_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X17 a_1003_n900# a_803_n964# a_745_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X18 a_745_n900# a_545_n964# a_487_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X19 a_487_n900# a_287_n964# a_229_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X20 a_1777_n900# a_1577_n964# a_1519_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
X21 a_2035_n900# a_1835_n964# a_1777_n900# w_n3067_n1197# sky130_fd_pr__pfet_g5v0d10v5 ad=1.305 pd=9.29 as=1.305 ps=9.29 w=9 l=1
C0 w_n3067_n1197# a_287_n964# 0.307639f
C1 a_n2867_n900# a_n2609_n900# 0.492143f
C2 a_n287_n900# a_n545_n900# 0.492143f
C3 a_n229_n964# a_n29_n900# 0.197777f
C4 a_n2809_n964# a_n2609_n900# 0.197777f
C5 a_2035_n900# a_2293_n900# 0.492143f
C6 a_n745_n964# a_n545_n900# 0.197777f
C7 a_1777_n900# a_1835_n964# 0.197777f
C8 a_229_n900# a_29_n964# 0.197777f
C9 a_n1003_n964# a_n803_n900# 0.197777f
C10 a_n1777_n964# a_n1835_n900# 0.197777f
C11 a_545_n964# w_n3067_n1197# 0.307639f
C12 a_2293_n900# a_2351_n964# 0.197777f
C13 w_n3067_n1197# a_2351_n964# 0.307639f
C14 a_n1519_n964# a_n1577_n900# 0.197777f
C15 a_1061_n964# a_1003_n900# 0.197777f
C16 a_229_n900# a_487_n900# 0.492143f
C17 a_n2351_n900# a_n2609_n900# 0.492143f
C18 a_1577_n964# w_n3067_n1197# 0.307639f
C19 a_n1003_n964# w_n3067_n1197# 0.307639f
C20 a_229_n900# a_287_n964# 0.197777f
C21 a_1319_n964# w_n3067_n1197# 0.307639f
C22 a_1061_n964# w_n3067_n1197# 0.307639f
C23 a_n29_n900# a_29_n964# 0.197777f
C24 a_n1519_n964# a_n1319_n900# 0.197777f
C25 w_n3067_n1197# a_n1261_n964# 0.307639f
C26 a_2093_n964# a_2293_n900# 0.197777f
C27 a_2093_n964# w_n3067_n1197# 0.307639f
C28 a_n2867_n900# a_n2809_n964# 0.197777f
C29 a_1261_n900# a_1003_n900# 0.492143f
C30 a_2035_n900# a_2093_n964# 0.197777f
C31 a_n2035_n964# a_n1835_n900# 0.197777f
C32 a_n803_n900# a_n1061_n900# 0.492143f
C33 a_2035_n900# a_1777_n900# 0.492143f
C34 a_n229_n964# a_n287_n900# 0.197777f
C35 a_n2351_n900# a_n2293_n964# 0.197777f
C36 a_n229_n964# w_n3067_n1197# 0.307639f
C37 a_n2093_n900# a_n1835_n900# 0.492143f
C38 a_n29_n900# a_n287_n900# 0.492143f
C39 a_n2293_n964# a_n2093_n900# 0.197777f
C40 a_1519_n900# a_1577_n964# 0.197777f
C41 a_n2351_n900# a_n2551_n964# 0.197777f
C42 a_745_n900# a_1003_n900# 0.492143f
C43 a_487_n900# a_745_n900# 0.492143f
C44 a_n2293_n964# w_n3067_n1197# 0.307639f
C45 a_1519_n900# a_1319_n964# 0.197777f
C46 a_2551_n900# a_2809_n900# 0.492143f
C47 a_n1319_n900# a_n1577_n900# 0.492143f
C48 a_n1777_n964# w_n3067_n1197# 0.307639f
C49 a_1577_n964# a_1777_n900# 0.197777f
C50 w_n3067_n1197# a_n2551_n964# 0.307639f
C51 a_1519_n900# a_1777_n900# 0.492143f
C52 a_n487_n964# a_n287_n900# 0.197777f
C53 a_745_n900# a_803_n964# 0.197777f
C54 a_n2867_n900# w_n3067_n1197# 0.529871f
C55 a_n1577_n900# a_n1835_n900# 0.492143f
C56 w_n3067_n1197# a_1835_n964# 0.307639f
C57 a_2035_n900# a_1835_n964# 0.197777f
C58 w_n3067_n1197# a_n2809_n964# 0.34286f
C59 a_n487_n964# w_n3067_n1197# 0.307639f
C60 a_2609_n964# a_2809_n900# 0.197777f
C61 a_n1319_n900# a_n1261_n964# 0.197777f
C62 a_2609_n964# a_2551_n900# 0.197777f
C63 a_29_n964# w_n3067_n1197# 0.307639f
C64 a_1519_n900# a_1261_n900# 0.492143f
C65 a_745_n900# a_545_n964# 0.197777f
C66 a_n487_n964# a_n545_n900# 0.197777f
C67 a_1261_n900# a_1319_n964# 0.197777f
C68 a_1261_n900# a_1061_n964# 0.197777f
C69 a_n1777_n964# a_n1577_n900# 0.197777f
C70 a_n745_n964# a_n803_n900# 0.197777f
C71 a_n1003_n964# a_n1061_n900# 0.197777f
C72 w_n3067_n1197# a_2809_n900# 0.529871f
C73 a_2551_n900# a_2293_n900# 0.492143f
C74 a_803_n964# a_1003_n900# 0.197777f
C75 a_n2093_n900# a_n2035_n964# 0.197777f
C76 a_487_n900# a_287_n964# 0.197777f
C77 a_n1061_n900# a_n1261_n964# 0.197777f
C78 w_n3067_n1197# a_n2035_n964# 0.307639f
C79 a_229_n900# a_n29_n900# 0.492143f
C80 a_n2351_n900# a_n2093_n900# 0.492143f
C81 a_2551_n900# a_2351_n964# 0.197777f
C82 a_n803_n900# a_n545_n900# 0.492143f
C83 a_n1519_n964# w_n3067_n1197# 0.307639f
C84 a_n1319_n900# a_n1061_n900# 0.492143f
C85 a_2609_n964# w_n3067_n1197# 0.34286f
C86 a_487_n900# a_545_n964# 0.197777f
C87 a_n2551_n964# a_n2609_n900# 0.197777f
C88 w_n3067_n1197# a_803_n964# 0.307639f
C89 a_n745_n964# w_n3067_n1197# 0.307639f
C90 a_2809_n900# 0 0.442831f
C91 a_2551_n900# 0 0.253417f
C92 a_2293_n900# 0 0.253417f
C93 a_2035_n900# 0 0.253417f
C94 a_1777_n900# 0 0.253417f
C95 a_1519_n900# 0 0.253417f
C96 a_1261_n900# 0 0.253417f
C97 a_1003_n900# 0 0.253417f
C98 a_745_n900# 0 0.253417f
C99 a_487_n900# 0 0.253417f
C100 a_229_n900# 0 0.253417f
C101 a_n29_n900# 0 0.253417f
C102 a_n287_n900# 0 0.253417f
C103 a_n545_n900# 0 0.253417f
C104 a_n803_n900# 0 0.253417f
C105 a_n1061_n900# 0 0.253417f
C106 a_n1319_n900# 0 0.253417f
C107 a_n1577_n900# 0 0.253417f
C108 a_n1835_n900# 0 0.253417f
C109 a_n2093_n900# 0 0.253417f
C110 a_n2351_n900# 0 0.253417f
C111 a_n2609_n900# 0 0.253417f
C112 a_n2867_n900# 0 0.442831f
C113 a_2609_n964# 0 0.253452f
C114 a_2351_n964# 0 0.231023f
C115 a_2093_n964# 0 0.231023f
C116 a_1835_n964# 0 0.231023f
C117 a_1577_n964# 0 0.231023f
C118 a_1319_n964# 0 0.231023f
C119 a_1061_n964# 0 0.231023f
C120 a_803_n964# 0 0.231023f
C121 a_545_n964# 0 0.231023f
C122 a_287_n964# 0 0.231023f
C123 a_29_n964# 0 0.231023f
C124 a_n229_n964# 0 0.231023f
C125 a_n487_n964# 0 0.231023f
C126 a_n745_n964# 0 0.231023f
C127 a_n1003_n964# 0 0.231023f
C128 a_n1261_n964# 0 0.231023f
C129 a_n1519_n964# 0 0.231023f
C130 a_n1777_n964# 0 0.231023f
C131 a_n2035_n964# 0 0.231023f
C132 a_n2293_n964# 0 0.231023f
C133 a_n2551_n964# 0 0.231023f
C134 a_n2809_n964# 0 0.253452f
C135 w_n3067_n1197# 0 48.853f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_HG2LSW a_n100_n205# a_100_n150# a_n292_n372#
+ a_n158_n150#
X0 a_100_n150# a_n100_n205# a_n158_n150# a_n292_n372# sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=1
C0 a_100_n150# a_n292_n372# 0.189446f
C1 a_n158_n150# a_n292_n372# 0.189446f
C2 a_n100_n205# a_n292_n372# 0.603705f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_N64HU4 a_3235_n255# a_n1861_n200# a_n1803_n255#
+ a_n3827_n422# a_n2777_n200# a_n1345_n255# a_n2719_n255# a_3635_n200# a_2261_n200#
+ a_n1403_n200# a_3177_n200# a_n2319_n200# a_1861_n255# a_2777_n255# a_1403_n255#
+ a_n887_n255# a_n945_n200# a_945_n255# a_2319_n255# a_n487_n200# a_n429_n255# a_1803_n200#
+ a_487_n255# a_2719_n200# a_1345_n200# a_n29_n200# a_n3693_n200# a_n2261_n255# a_n3635_n255#
+ a_887_n200# a_29_n255# a_n3177_n255# a_n3235_n200# a_429_n200#
X0 a_1345_n200# a_945_n255# a_887_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X1 a_n2319_n200# a_n2719_n255# a_n2777_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X2 a_n2777_n200# a_n3177_n255# a_n3235_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X3 a_2261_n200# a_1861_n255# a_1803_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X4 a_n945_n200# a_n1345_n255# a_n1403_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X5 a_3635_n200# a_3235_n255# a_3177_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X6 a_429_n200# a_29_n255# a_n29_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X7 a_1803_n200# a_1403_n255# a_1345_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X8 a_887_n200# a_487_n255# a_429_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X9 a_3177_n200# a_2777_n255# a_2719_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X10 a_n3235_n200# a_n3635_n255# a_n3693_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X11 a_n487_n200# a_n887_n255# a_n945_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X12 a_n1403_n200# a_n1803_n255# a_n1861_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X13 a_2719_n200# a_2319_n255# a_2261_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X14 a_n1861_n200# a_n2261_n255# a_n2319_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X15 a_n29_n200# a_n429_n255# a_n487_n200# a_n3827_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
C0 a_3635_n200# a_n3827_n422# 0.256295f
C1 a_3177_n200# a_n3827_n422# 0.114065f
C2 a_2719_n200# a_n3827_n422# 0.114065f
C3 a_2261_n200# a_n3827_n422# 0.114065f
C4 a_1803_n200# a_n3827_n422# 0.114065f
C5 a_1345_n200# a_n3827_n422# 0.114065f
C6 a_887_n200# a_n3827_n422# 0.114065f
C7 a_429_n200# a_n3827_n422# 0.114065f
C8 a_n29_n200# a_n3827_n422# 0.114065f
C9 a_n487_n200# a_n3827_n422# 0.114065f
C10 a_n945_n200# a_n3827_n422# 0.114065f
C11 a_n1403_n200# a_n3827_n422# 0.114065f
C12 a_n1861_n200# a_n3827_n422# 0.114065f
C13 a_n2319_n200# a_n3827_n422# 0.114065f
C14 a_n2777_n200# a_n3827_n422# 0.114065f
C15 a_n3235_n200# a_n3827_n422# 0.114065f
C16 a_n3693_n200# a_n3827_n422# 0.256295f
C17 a_3235_n255# a_n3827_n422# 0.994274f
C18 a_2777_n255# a_n3827_n422# 0.946497f
C19 a_2319_n255# a_n3827_n422# 0.946497f
C20 a_1861_n255# a_n3827_n422# 0.946497f
C21 a_1403_n255# a_n3827_n422# 0.946497f
C22 a_945_n255# a_n3827_n422# 0.946497f
C23 a_487_n255# a_n3827_n422# 0.946497f
C24 a_29_n255# a_n3827_n422# 0.946497f
C25 a_n429_n255# a_n3827_n422# 0.946497f
C26 a_n887_n255# a_n3827_n422# 0.946497f
C27 a_n1345_n255# a_n3827_n422# 0.946497f
C28 a_n1803_n255# a_n3827_n422# 0.946497f
C29 a_n2261_n255# a_n3827_n422# 0.946497f
C30 a_n2719_n255# a_n3827_n422# 0.946497f
C31 a_n3177_n255# a_n3827_n422# 0.946497f
C32 a_n3635_n255# a_n3827_n422# 0.994274f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_RMXH5H a_803_n255# a_1261_n200# a_n1319_n200#
+ a_n287_n200# a_n229_n255# a_n1061_n200# a_287_n255# a_n1003_n255# a_745_n200# a_1319_n255#
+ a_n1711_n422# a_1061_n255# a_229_n200# a_n1577_n200# a_n1519_n255# a_n487_n255#
+ a_n545_n200# a_n1261_n255# a_545_n255# a_1003_n200# a_487_n200# a_n29_n200# a_29_n255#
+ a_n745_n255# a_n803_n200# a_1519_n200#
X0 a_487_n200# a_287_n255# a_229_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X1 a_1261_n200# a_1061_n255# a_1003_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X2 a_n29_n200# a_n229_n255# a_n287_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X3 a_229_n200# a_29_n255# a_n29_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X4 a_n1319_n200# a_n1519_n255# a_n1577_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X5 a_n545_n200# a_n745_n255# a_n803_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X6 a_n803_n200# a_n1003_n255# a_n1061_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X7 a_n287_n200# a_n487_n255# a_n545_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X8 a_1519_n200# a_1319_n255# a_1261_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X9 a_n1061_n200# a_n1261_n255# a_n1319_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X10 a_745_n200# a_545_n255# a_487_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
X11 a_1003_n200# a_803_n255# a_745_n200# a_n1711_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=1
C0 a_1261_n200# a_1003_n200# 0.110175f
C1 a_487_n200# a_229_n200# 0.110175f
C2 a_n1577_n200# a_n1319_n200# 0.110175f
C3 a_n29_n200# a_229_n200# 0.110175f
C4 a_n1319_n200# a_n1061_n200# 0.110175f
C5 a_n545_n200# a_n803_n200# 0.110175f
C6 a_487_n200# a_745_n200# 0.110175f
C7 a_n545_n200# a_n287_n200# 0.110175f
C8 a_n1061_n200# a_n803_n200# 0.110175f
C9 a_1519_n200# a_1261_n200# 0.110175f
C10 a_n287_n200# a_n29_n200# 0.110175f
C11 a_745_n200# a_1003_n200# 0.110175f
C12 a_1519_n200# a_n1711_n422# 0.241444f
C13 a_n1577_n200# a_n1711_n422# 0.241444f
C14 a_1319_n255# a_n1711_n422# 0.55256f
C15 a_1061_n255# a_n1711_n422# 0.498389f
C16 a_803_n255# a_n1711_n422# 0.498389f
C17 a_545_n255# a_n1711_n422# 0.498389f
C18 a_287_n255# a_n1711_n422# 0.498389f
C19 a_29_n255# a_n1711_n422# 0.498389f
C20 a_n229_n255# a_n1711_n422# 0.498389f
C21 a_n487_n255# a_n1711_n422# 0.498389f
C22 a_n745_n255# a_n1711_n422# 0.498389f
C23 a_n1003_n255# a_n1711_n422# 0.498389f
C24 a_n1261_n255# a_n1711_n422# 0.498389f
C25 a_n1519_n255# a_n1711_n422# 0.55256f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_TT9EEV a_n932_n420# a_1648_n420# a_n1648_n484#
+ a_1390_n420# a_n1390_n484# a_n616_n484# a_n1448_n420# a_674_n484# a_n1190_n420#
+ w_n1906_n717# a_n416_n420# a_874_n420# a_158_n484# a_358_n420# a_n874_n484# a_n1706_n420#
+ a_932_n484# a_100_n420# a_n674_n420# a_1132_n420# a_n358_n484# a_n1132_n484# a_416_n484#
+ a_n158_n420# a_n100_n484# a_616_n420# a_1448_n484# a_1190_n484#
X0 a_n416_n420# a_n616_n484# a_n674_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X1 a_n158_n420# a_n358_n484# a_n416_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X2 a_n1448_n420# a_n1648_n484# a_n1706_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=1.218 ps=8.98 w=4.2 l=1
X3 a_n1190_n420# a_n1390_n484# a_n1448_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X4 a_n674_n420# a_n874_n484# a_n932_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X5 a_n932_n420# a_n1132_n484# a_n1190_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X6 a_358_n420# a_158_n484# a_100_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X7 a_616_n420# a_416_n484# a_358_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X8 a_1648_n420# a_1448_n484# a_1390_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=1.218 pd=8.98 as=0.609 ps=4.49 w=4.2 l=1
X9 a_1132_n420# a_932_n484# a_874_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X10 a_874_n420# a_674_n484# a_616_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X11 a_1390_n420# a_1190_n484# a_1132_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
X12 a_100_n420# a_n100_n484# a_n158_n420# w_n1906_n717# sky130_fd_pr__pfet_g5v0d10v5 ad=0.609 pd=4.49 as=0.609 ps=4.49 w=4.2 l=1
C0 w_n1906_n717# a_n1648_n484# 0.34286f
C1 a_n674_n420# a_n416_n420# 0.230222f
C2 a_1390_n420# a_1648_n420# 0.230222f
C3 w_n1906_n717# a_n358_n484# 0.307639f
C4 a_358_n420# a_100_n420# 0.230222f
C5 a_n158_n420# a_100_n420# 0.230222f
C6 w_n1906_n717# a_n874_n484# 0.307639f
C7 w_n1906_n717# a_n100_n484# 0.307639f
C8 w_n1906_n717# a_932_n484# 0.307639f
C9 a_n1190_n420# a_n932_n420# 0.230222f
C10 a_n158_n420# a_n416_n420# 0.230222f
C11 w_n1906_n717# a_n1706_n420# 0.260562f
C12 a_1390_n420# a_1132_n420# 0.230222f
C13 w_n1906_n717# a_158_n484# 0.307639f
C14 a_n1190_n420# a_n1448_n420# 0.230222f
C15 w_n1906_n717# a_1448_n484# 0.34286f
C16 a_n932_n420# a_n674_n420# 0.230222f
C17 a_n1706_n420# a_n1448_n420# 0.230222f
C18 a_n1390_n484# w_n1906_n717# 0.307639f
C19 w_n1906_n717# a_674_n484# 0.307639f
C20 w_n1906_n717# a_n1132_n484# 0.307639f
C21 a_874_n420# a_1132_n420# 0.230222f
C22 w_n1906_n717# a_1648_n420# 0.260562f
C23 w_n1906_n717# a_416_n484# 0.307639f
C24 a_616_n420# a_358_n420# 0.230222f
C25 a_874_n420# a_616_n420# 0.230222f
C26 w_n1906_n717# a_n616_n484# 0.307639f
C27 a_1190_n484# w_n1906_n717# 0.307639f
C28 a_1648_n420# 0 0.211168f
C29 a_1390_n420# 0 0.122326f
C30 a_1132_n420# 0 0.122326f
C31 a_874_n420# 0 0.122326f
C32 a_616_n420# 0 0.122326f
C33 a_358_n420# 0 0.122326f
C34 a_100_n420# 0 0.122326f
C35 a_n158_n420# 0 0.122326f
C36 a_n416_n420# 0 0.122326f
C37 a_n674_n420# 0 0.122326f
C38 a_n932_n420# 0 0.122326f
C39 a_n1190_n420# 0 0.122326f
C40 a_n1448_n420# 0 0.122326f
C41 a_n1706_n420# 0 0.211168f
C42 a_1448_n484# 0 0.234278f
C43 a_1190_n484# 0 0.211849f
C44 a_932_n484# 0 0.211849f
C45 a_674_n484# 0 0.211849f
C46 a_416_n484# 0 0.211849f
C47 a_158_n484# 0 0.211849f
C48 a_n100_n484# 0 0.211849f
C49 a_n358_n484# 0 0.211849f
C50 a_n616_n484# 0 0.211849f
C51 a_n874_n484# 0 0.211849f
C52 a_n1132_n484# 0 0.211849f
C53 a_n1390_n484# 0 0.211849f
C54 a_n1648_n484# 0 0.234278f
C55 w_n1906_n717# 0 19.199598f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_BH2H9S a_n229_n1664# a_1061_n1664# a_n1835_n1600#
+ a_n2351_n1600# a_n1261_n1664# a_n1061_n1600# a_1319_n1664# a_1261_n1600# a_287_n1664#
+ a_n2035_n1664# a_2035_n1600# a_n1319_n1600# a_n1519_n1664# a_1519_n1600# a_487_n1600#
+ a_545_n1664# a_29_n1664# a_n487_n1664# a_n287_n1600# w_n2551_n1897# a_745_n1600#
+ a_2093_n1664# a_1577_n1664# a_803_n1664# a_n745_n1664# a_n1003_n1664# a_1003_n1600#
+ a_n545_n1600# a_n2293_n1664# a_n2093_n1600# a_n1777_n1664# a_2293_n1600# a_n1577_n1600#
+ a_1777_n1600# a_n29_n1600# a_1835_n1664# a_229_n1600# a_n803_n1600#
X0 a_n287_n1600# a_n487_n1664# a_n545_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X1 a_n1577_n1600# a_n1777_n1664# a_n1835_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X2 a_n29_n1600# a_n229_n1664# a_n287_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X3 a_2035_n1600# a_1835_n1664# a_1777_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X4 a_n1319_n1600# a_n1519_n1664# a_n1577_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X5 a_n2093_n1600# a_n2293_n1664# a_n2351_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=1
X6 a_745_n1600# a_545_n1664# a_487_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X7 a_n1835_n1600# a_n2035_n1664# a_n2093_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X8 a_1261_n1600# a_1061_n1664# a_1003_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X9 a_n545_n1600# a_n745_n1664# a_n803_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X10 a_229_n1600# a_29_n1664# a_n29_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X11 a_1003_n1600# a_803_n1664# a_745_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X12 a_n1061_n1600# a_n1261_n1664# a_n1319_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X13 a_n803_n1600# a_n1003_n1664# a_n1061_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X14 a_1777_n1600# a_1577_n1664# a_1519_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X15 a_1519_n1600# a_1319_n1664# a_1261_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X16 a_487_n1600# a_287_n1664# a_229_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=1
X17 a_2293_n1600# a_2093_n1664# a_2035_n1600# w_n2551_n1897# sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=1
C0 a_1519_n1600# a_1777_n1600# 0.874111f
C1 a_229_n1600# a_n29_n1600# 0.874111f
C2 a_229_n1600# a_29_n1664# 0.347373f
C3 a_n1319_n1600# a_n1061_n1600# 0.874111f
C4 a_n1061_n1600# a_n1003_n1664# 0.347373f
C5 a_n2351_n1600# a_n2293_n1664# 0.347373f
C6 a_n1319_n1600# a_n1577_n1600# 0.874111f
C7 w_n2551_n1897# a_n1261_n1664# 0.307639f
C8 w_n2551_n1897# a_n1519_n1664# 0.307639f
C9 a_487_n1600# a_745_n1600# 0.874111f
C10 a_2035_n1600# a_2293_n1600# 0.874111f
C11 w_n2551_n1897# a_803_n1664# 0.307639f
C12 w_n2551_n1897# a_2293_n1600# 0.922614f
C13 a_n2093_n1600# a_n2351_n1600# 0.874111f
C14 w_n2551_n1897# a_n745_n1664# 0.307639f
C15 a_n545_n1600# a_n745_n1664# 0.347373f
C16 a_n803_n1600# a_n745_n1664# 0.347373f
C17 a_1261_n1600# a_1061_n1664# 0.347373f
C18 a_1319_n1664# w_n2551_n1897# 0.307639f
C19 a_n2093_n1600# a_n1835_n1600# 0.874111f
C20 a_2093_n1664# a_2035_n1600# 0.347373f
C21 w_n2551_n1897# a_2093_n1664# 0.34286f
C22 a_n803_n1600# a_n1061_n1600# 0.874111f
C23 a_1003_n1600# a_1061_n1664# 0.347373f
C24 a_1003_n1600# a_1261_n1600# 0.874111f
C25 a_n287_n1600# a_n229_n1664# 0.347373f
C26 a_1519_n1600# a_1577_n1664# 0.347373f
C27 w_n2551_n1897# a_n1777_n1664# 0.307639f
C28 w_n2551_n1897# a_n229_n1664# 0.307639f
C29 w_n2551_n1897# a_n2035_n1664# 0.307639f
C30 a_2035_n1600# a_1777_n1600# 0.874111f
C31 a_1835_n1664# a_1777_n1600# 0.347373f
C32 w_n2551_n1897# a_n1003_n1664# 0.307639f
C33 a_n29_n1600# a_29_n1664# 0.347373f
C34 a_n803_n1600# a_n1003_n1664# 0.347373f
C35 a_1777_n1600# a_1577_n1664# 0.347373f
C36 a_545_n1664# a_745_n1600# 0.347373f
C37 a_n2093_n1600# a_n2035_n1664# 0.347373f
C38 a_2035_n1600# a_1835_n1664# 0.347373f
C39 a_1003_n1600# a_745_n1600# 0.874111f
C40 a_1319_n1664# a_1261_n1600# 0.347373f
C41 a_1003_n1600# a_803_n1664# 0.347373f
C42 w_n2551_n1897# a_1835_n1664# 0.307639f
C43 a_n287_n1600# a_n545_n1600# 0.874111f
C44 a_1261_n1600# a_1519_n1600# 0.874111f
C45 a_n803_n1600# a_n545_n1600# 0.874111f
C46 a_487_n1600# a_229_n1600# 0.874111f
C47 w_n2551_n1897# a_1577_n1664# 0.307639f
C48 w_n2551_n1897# a_n2293_n1664# 0.34286f
C49 a_n229_n1664# a_n29_n1600# 0.347373f
C50 a_803_n1664# a_745_n1600# 0.347373f
C51 a_n1835_n1600# a_n1577_n1600# 0.874111f
C52 a_n287_n1600# a_n487_n1664# 0.347373f
C53 w_n2551_n1897# a_n487_n1664# 0.307639f
C54 a_n1061_n1600# a_n1261_n1664# 0.347373f
C55 a_n545_n1600# a_n487_n1664# 0.347373f
C56 a_n1835_n1600# a_n1777_n1664# 0.347373f
C57 a_n1519_n1664# a_n1577_n1600# 0.347373f
C58 a_n2035_n1664# a_n1835_n1600# 0.347373f
C59 a_487_n1600# a_545_n1664# 0.347373f
C60 a_n2093_n1600# a_n2293_n1664# 0.347373f
C61 w_n2551_n1897# a_545_n1664# 0.307639f
C62 a_2093_n1664# a_2293_n1600# 0.347373f
C63 a_1319_n1664# a_1519_n1600# 0.347373f
C64 w_n2551_n1897# a_1061_n1664# 0.307639f
C65 a_487_n1600# a_287_n1664# 0.347373f
C66 a_n1319_n1600# a_n1261_n1664# 0.347373f
C67 a_n1519_n1664# a_n1319_n1600# 0.347373f
C68 w_n2551_n1897# a_287_n1664# 0.307639f
C69 a_n287_n1600# a_n29_n1600# 0.874111f
C70 a_229_n1600# a_287_n1664# 0.347373f
C71 w_n2551_n1897# a_29_n1664# 0.307639f
C72 w_n2551_n1897# a_n2351_n1600# 0.922614f
C73 a_n1777_n1664# a_n1577_n1600# 0.347373f
C74 a_2293_n1600# 0 0.780672f
C75 a_2035_n1600# 0 0.44459f
C76 a_1777_n1600# 0 0.44459f
C77 a_1519_n1600# 0 0.44459f
C78 a_1261_n1600# 0 0.44459f
C79 a_1003_n1600# 0 0.44459f
C80 a_745_n1600# 0 0.44459f
C81 a_487_n1600# 0 0.44459f
C82 a_229_n1600# 0 0.44459f
C83 a_n29_n1600# 0 0.44459f
C84 a_n287_n1600# 0 0.44459f
C85 a_n545_n1600# 0 0.44459f
C86 a_n803_n1600# 0 0.44459f
C87 a_n1061_n1600# 0 0.44459f
C88 a_n1319_n1600# 0 0.44459f
C89 a_n1577_n1600# 0 0.44459f
C90 a_n1835_n1600# 0 0.44459f
C91 a_n2093_n1600# 0 0.44459f
C92 a_n2351_n1600# 0 0.780672f
C93 a_2093_n1664# 0 0.253452f
C94 a_1835_n1664# 0 0.231023f
C95 a_1577_n1664# 0 0.231023f
C96 a_1319_n1664# 0 0.231023f
C97 a_1061_n1664# 0 0.231023f
C98 a_803_n1664# 0 0.231023f
C99 a_545_n1664# 0 0.231023f
C100 a_287_n1664# 0 0.231023f
C101 a_29_n1664# 0 0.231023f
C102 a_n229_n1664# 0 0.231023f
C103 a_n487_n1664# 0 0.231023f
C104 a_n745_n1664# 0 0.231023f
C105 a_n1003_n1664# 0 0.231023f
C106 a_n1261_n1664# 0 0.231023f
C107 a_n1519_n1664# 0 0.231023f
C108 a_n1777_n1664# 0 0.231023f
C109 a_n2035_n1664# 0 0.231023f
C110 a_n2293_n1664# 0 0.253452f
C111 w_n2551_n1897# 0 62.9271f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U a_n1861_n200# a_n1803_n255# a_n3369_n422#
+ a_n2777_n200# a_n1345_n255# a_n2719_n255# a_2261_n200# a_n1403_n200# a_3177_n200#
+ a_n2319_n200# a_1861_n255# a_2777_n255# a_1403_n255# a_n887_n255# a_n945_n200# a_945_n255#
+ a_2319_n255# a_n487_n200# a_n429_n255# a_1803_n200# a_487_n255# a_2719_n200# a_1345_n200#
+ a_n29_n200# a_n2261_n255# a_887_n200# a_29_n255# a_n3177_n255# a_n3235_n200# a_429_n200#
X0 a_1345_n200# a_945_n255# a_887_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X1 a_n2319_n200# a_n2719_n255# a_n2777_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X2 a_n2777_n200# a_n3177_n255# a_n3235_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=2
X3 a_2261_n200# a_1861_n255# a_1803_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X4 a_n945_n200# a_n1345_n255# a_n1403_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X5 a_429_n200# a_29_n255# a_n29_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X6 a_1803_n200# a_1403_n255# a_1345_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X7 a_887_n200# a_487_n255# a_429_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X8 a_3177_n200# a_2777_n255# a_2719_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=2
X9 a_n487_n200# a_n887_n255# a_n945_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X10 a_n1403_n200# a_n1803_n255# a_n1861_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X11 a_2719_n200# a_2319_n255# a_2261_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X12 a_n1861_n200# a_n2261_n255# a_n2319_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
X13 a_n29_n200# a_n429_n255# a_n487_n200# a_n3369_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=2
C0 a_3177_n200# a_n3369_n422# 0.256295f
C1 a_2719_n200# a_n3369_n422# 0.114065f
C2 a_2261_n200# a_n3369_n422# 0.114065f
C3 a_1803_n200# a_n3369_n422# 0.114065f
C4 a_1345_n200# a_n3369_n422# 0.114065f
C5 a_887_n200# a_n3369_n422# 0.114065f
C6 a_429_n200# a_n3369_n422# 0.114065f
C7 a_n29_n200# a_n3369_n422# 0.114065f
C8 a_n487_n200# a_n3369_n422# 0.114065f
C9 a_n945_n200# a_n3369_n422# 0.114065f
C10 a_n1403_n200# a_n3369_n422# 0.114065f
C11 a_n1861_n200# a_n3369_n422# 0.114065f
C12 a_n2319_n200# a_n3369_n422# 0.114065f
C13 a_n2777_n200# a_n3369_n422# 0.114065f
C14 a_n3235_n200# a_n3369_n422# 0.256295f
C15 a_2777_n255# a_n3369_n422# 0.994274f
C16 a_2319_n255# a_n3369_n422# 0.946497f
C17 a_1861_n255# a_n3369_n422# 0.946497f
C18 a_1403_n255# a_n3369_n422# 0.946497f
C19 a_945_n255# a_n3369_n422# 0.946497f
C20 a_487_n255# a_n3369_n422# 0.946497f
C21 a_29_n255# a_n3369_n422# 0.946497f
C22 a_n429_n255# a_n3369_n422# 0.946497f
C23 a_n887_n255# a_n3369_n422# 0.946497f
C24 a_n1345_n255# a_n3369_n422# 0.946497f
C25 a_n1803_n255# a_n3369_n422# 0.946497f
C26 a_n2261_n255# a_n3369_n422# 0.946497f
C27 a_n2719_n255# a_n3369_n422# 0.946497f
C28 a_n3177_n255# a_n3369_n422# 0.994274f
.ends

.subckt sky130_td_ip__opamp_hp avdd vout ibias vinn vinp dvdd dvss ena avss
Xsky130_fd_pr__pfet_g5v0d10v5_W75H7K_0 m1_180_3630# avdd m1_n1154_3624# m1_n1154_3624#
+ avdd m1_180_3630# avdd m1_n1154_3624# m1_n1154_3624# m1_n1154_3624# m1_n1154_3624#
+ m1_806_3964# m1_n1154_3624# m1_n1154_3624# m1_806_3964# m1_180_3630# avdd avdd m1_n1154_3624#
+ m1_n1154_3624# avdd m1_180_3630# m1_806_3964# avdd m1_n1154_3624# m1_n1154_3624#
+ m1_n1154_3624# avdd m1_806_3964# m1_180_3630# m1_n1154_3624# avdd avdd m1_n1154_3624#
+ m1_n1154_3624# avdd m1_806_3964# m1_n1154_3624# avdd m1_n1154_3624# m1_n1154_3624#
+ m1_180_3630# m1_n1154_3624# m1_n1154_3624# avdd m1_n1154_3624# m1_806_3964# avdd
+ m1_n1154_3624# m1_180_3630# avdd m1_n1154_3624# m1_n1154_3624# avdd m1_180_3630#
+ m1_n1154_3624# m1_n1154_3624# m1_n1154_3624# m1_180_3630# m1_n1154_3624# avdd m1_806_3964#
+ avdd m1_n1154_3624# m1_806_3964# m1_n1154_3624# m1_180_3630# avdd m1_806_3964# avdd
+ avdd m1_n1154_3624# m1_n1154_3624# m1_n1154_3624# avdd m1_n1154_3624# m1_n1154_3624#
+ avdd sky130_fd_pr__pfet_g5v0d10v5_W75H7K
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_15 avdd avdd m1_n1846_3922# m1_n3561_8311# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_16 m1_n1154_3624# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_WKXP7K_0 m1_806_3964# m1_n592_3104# avdd m1_790_6356#
+ m1_790_6356# m1_180_3630# m1_n592_3104# m1_790_6356# m1_790_6356# m1_790_6356# m1_790_6356#
+ m1_806_3964# m1_790_6356# m1_790_6356# m1_180_3630# m1_180_3630# m1_n1154_3624#
+ m1_n1154_3624# m1_790_6356# m1_790_6356# m1_n592_3104# m1_806_3964# m1_806_3964#
+ m1_n1154_3624# m1_790_6356# m1_790_6356# m1_790_6356# m1_n592_3104# avdd m1_806_3964#
+ m1_790_6356# m1_n592_3104# m1_n1154_3624# m1_790_6356# m1_790_6356# m1_n592_3104#
+ m1_806_3964# avdd m1_n592_3104# m1_790_6356# m1_790_6356# m1_180_3630# m1_790_6356#
+ m1_790_6356# m1_n1154_3624# m1_790_6356# avdd avdd avdd m1_180_3630# m1_n1154_3624#
+ m1_790_6356# m1_180_3630# m1_n1154_3624# m1_790_6356# m1_790_6356# m1_n592_3104#
+ m1_806_3964# m1_790_6356# m1_790_6356# m1_790_6356# m1_806_3964# m1_790_6356# m1_n592_3104#
+ m1_806_3964# m1_n592_3104# m1_790_6356# m1_180_3630# m1_790_6356# m1_180_3630# m1_n1154_3624#
+ m1_180_3630# m1_n1154_3624# m1_790_6356# m1_790_6356# avdd m1_790_6356# m1_n1154_3624#
+ m1_790_6356# avdd m1_790_6356# m1_790_6356# sky130_fd_pr__pfet_g5v0d10v5_WKXP7K
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_17 m1_n1846_3922# avdd m1_n3264_4838# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_01v8_6H2JYD_0 dvss m1_n9267_3854# m1_n8442_3847# dvss sky130_fd_pr__nfet_01v8_6H2JYD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_0 ibias avss m1_n3955_n943# m1_n3750_n668# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_HQ4STX_0 avdd m1_790_6356# m1_790_6356# avdd sky130_fd_pr__pfet_g5v0d10v5_HQ4STX
Xsky130_fd_pr__nfet_01v8_6H2JYD_1 dvss ena m1_n9267_3854# dvss sky130_fd_pr__nfet_01v8_6H2JYD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_1 m1_n4685_n1863# avss m1_n4698_n3450# m1_n3750_n668#
+ sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_2 m1_n1846_3922# avss avss m1_n3264_4838# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_YJ3VXJ_0 m1_n8442_3847# m1_n3264_4838# avss avss avss
+ avss m1_n3264_4838# avss avss m1_n3667_4379# m1_n9267_3854# avss m1_n9267_3854#
+ m1_n8442_3847# sky130_fd_pr__nfet_g5v0d10v5_YJ3VXJ
Xsky130_fd_pr__nfet_g5v0d10v5_UKVZ7J_0 net29 avss net12 m1_n4692_n1074# avss m1_n4692_n1074#
+ m1_n4692_n1074# m1_n4692_n1074# avss avss net12 m1_n4692_n1074# m1_n4692_n1074#
+ avss m1_n4692_n1074# m1_n4692_n1074# avss avss net12 avss m1_n4692_n1074# net12
+ avss net12 m1_n4692_n1074# m1_n4692_n1074# avss m1_n4692_n1074# m1_n4692_n1074#
+ avss net29 avss net12 m1_n4692_n1074# net28 m1_n4692_n1074# m1_n4692_n1074# avss
+ net12 m1_n4692_n1074# avss m1_n4692_n1074# avss m1_n4692_n1074# m1_n4692_n1074#
+ net12 m1_n4692_n1074# net28 m1_n4692_n1074# avss avss net12 m1_n4692_n1074# m1_n4692_n1074#
+ sky130_fd_pr__nfet_g5v0d10v5_UKVZ7J
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_3 m1_n4694_n312# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_USXRNR_0 avss m1_n4704_472# avss avss avss m1_n4694_n312#
+ m1_n1154_3624# m1_n4704_472# m1_n4704_472# m1_n4704_472# m1_16202_3432# m1_n1154_3624#
+ avss m1_16202_3432# m1_n4704_472# m1_n4694_n312# avss m1_n4704_472# m1_n592_3104#
+ m1_n4694_n312# m1_n4704_472# m1_n4694_n312# m1_n1154_3624# m1_n4704_472# m1_n592_3104#
+ avss m1_n4704_472# avss sky130_fd_pr__nfet_g5v0d10v5_USXRNR
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_0 avdd avdd m1_n1846_3922# m1_806_3964# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_4 m1_n4704_472# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_1 m1_n3080_8896# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_5 vb3 avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_2 avdd avdd m1_n1846_3922# m1_779_5148# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_6 m1_n4692_n1074# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_AUMBFF_0 m1_n592_3104# m1_n592_3104# avdd vout avdd
+ vout avdd m1_n592_3104# m1_n592_3104# m1_n592_3104# vout m1_n592_3104# m1_n592_3104#
+ m1_n592_3104# m1_n592_3104# vout m1_n592_3104# m1_n592_3104# m1_n592_3104# avdd
+ avdd avdd avdd m1_n592_3104# m1_n592_3104# avdd vout avdd vout m1_n592_3104# m1_n592_3104#
+ vout avdd m1_n592_3104# vout avdd avdd avdd m1_n592_3104# avdd avdd m1_n592_3104#
+ vout vout m1_n592_3104# m1_n592_3104# vout avdd m1_n592_3104# m1_n592_3104# avdd
+ m1_n592_3104# m1_n592_3104# vout m1_n592_3104# avdd vout avdd m1_n592_3104# m1_n592_3104#
+ vout avdd m1_n592_3104# avdd m1_n592_3104# m1_n592_3104# m1_n592_3104# vout avdd
+ vout sky130_fd_pr__pfet_g5v0d10v5_AUMBFF
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_3 m1_n3777_8065# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_7 m1_n4685_n1863# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QL2RRT_0 vinn vinn m1_n5902_n1890# vinp m1_n5902_n1890#
+ m1_n2158_9110# vinp m1_n2158_9110# vinp vinn m1_n2158_9110# avdd vinn m1_n2158_9110#
+ vinn avdd vinn vinp m1_n5904_n2678# avdd vinn avdd m1_n2158_9110# m1_n2158_9110#
+ vinp m1_n5902_n1890# m1_n2158_9110# vinn m1_n5902_n1890# vinp m1_n5904_n2678# m1_n2158_9110#
+ m1_n2158_9110# vinp m1_n5904_n2678# vinn vinp vinp vinp m1_n5904_n2678# m1_n5902_n1890#
+ m1_n2158_9110# vinn m1_n5904_n2678# vinn m1_n5904_n2678# avdd vinp m1_n2158_9110#
+ vinn m1_n2158_9110# m1_n5902_n1890# m1_n2158_9110# vinp sky130_fd_pr__pfet_g5v0d10v5_QL2RRT
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_4 m1_n4182_7627# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_8 m1_n4700_n2510# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QL2RRT_1 vinp vinp m1_n5904_n2678# vinn m1_n5904_n2678#
+ m1_n2158_9110# vinn m1_n2158_9110# vinn vinp m1_n2158_9110# avdd vinp m1_n2158_9110#
+ vinp avdd vinp vinn m1_n5902_n1890# avdd vinp avdd m1_n2158_9110# m1_n2158_9110#
+ vinn m1_n5904_n2678# m1_n2158_9110# vinp m1_n5904_n2678# vinn m1_n5902_n1890# m1_n2158_9110#
+ m1_n2158_9110# vinn m1_n5902_n1890# vinp vinn vinn vinn m1_n5902_n1890# m1_n5904_n2678#
+ m1_n2158_9110# vinp m1_n5902_n1890# vinp m1_n5902_n1890# avdd vinn m1_n2158_9110#
+ vinp m1_n2158_9110# m1_n5904_n2678# m1_n2158_9110# vinn sky130_fd_pr__pfet_g5v0d10v5_QL2RRT
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_5 avdd avdd m1_n3667_4379# m1_n6000_2704# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_9 m1_n4698_n3450# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_7 avdd avdd m1_n1846_3922# m1_791_7588# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_6 avdd avdd m1_n1846_3922# m1_790_6356# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_8 m1_180_4838# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_01v8_U4BBJH_0 m1_n8442_3847# dvdd m1_n9267_3854# dvss dvdd sky130_fd_pr__pfet_01v8_U4BBJH
Xsky130_fd_pr__pfet_01v8_U4BBJH_1 m1_n9267_3854# dvdd ena dvss dvdd sky130_fd_pr__pfet_01v8_U4BBJH
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_9 m1_180_3630# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_QTY6KC_0 m1_18668_3467# m1_180_4838# m1_18668_3467#
+ avdd avdd avdd m1_18668_3467# avdd m1_18668_3467# avdd avdd m1_180_4838# m1_180_4838#
+ m1_18668_3467# m1_18668_3467# m1_18668_3467# m1_180_4838# avdd avdd m1_180_4838#
+ avdd avdd m1_18668_3467# m1_180_4838# m1_18668_3467# avdd sky130_fd_pr__pfet_g5v0d10v5_QTY6KC
Xsky130_fd_pr__nfet_g5v0d10v5_B3XH3Z_0 li_9924_630# avss m1_779_5148# avss net12 vb3
+ vb3 vb3 net29 avss li_9924_630# avss net12 m1_779_5148# vb3 avss net12 vb3 vb3 net12
+ net28 avss li_9924_630# vb3 vb3 li_9924_630# net12 m1_n4692_n1074# vb3 avss avss
+ vb3 vb3 net12 m1_779_5148# vb3 li_9924_630# avss vb3 li_9924_630# avss vb3 avss
+ li_9924_630# m1_n4692_n1074# vb3 vb3 net28 vb3 net12 vb3 vb3 li_9924_630# vb3 li_9924_630#
+ vb3 vb3 net12 net29 m1_n4692_n1074# vb3 vb3 sky130_fd_pr__nfet_g5v0d10v5_B3XH3Z
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_10 net12 avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QTY6H6_0 avdd m1_13086_11886# m1_13086_11886# avdd m1_13086_11886#
+ avdd m1_n3445_8429# avdd m1_13086_11886# avdd m1_13086_11886# avdd m1_13086_11886#
+ m1_n3445_8429# m1_n3445_8429# m1_13086_11886# m1_13086_11886# m1_13086_11886# m1_n3445_8429#
+ m1_n3208_8640# avdd m1_13086_11886# avdd avdd avdd avdd sky130_fd_pr__pfet_g5v0d10v5_QTY6H6
Xsky130_fd_pr__nfet_g5v0d10v5_U73S5M_0 vout vout m1_16202_3432# m1_16202_3432# m1_16202_3432#
+ avss avss vout avss m1_16202_3432# m1_16202_3432# avss vout vout avss m1_16202_3432#
+ m1_16202_3432# m1_16202_3432# m1_16202_3432# m1_16202_3432# m1_16202_3432# avss
+ avss m1_16202_3432# vout avss m1_16202_3432# vout vout avss m1_16202_3432# m1_16202_3432#
+ avss m1_16202_3432# avss avss vout vout m1_16202_3432# avss m1_16202_3432# m1_16202_3432#
+ vout m1_16202_3432# m1_16202_3432# m1_16202_3432# m1_16202_3432# m1_16202_3432#
+ m1_16202_3432# m1_16202_3432# avss vout m1_16202_3432# avss avss m1_16202_3432#
+ m1_16202_3432# m1_16202_3432# avss vout vout m1_16202_3432# avss m1_16202_3432#
+ vout avss avss vout avss avss sky130_fd_pr__nfet_g5v0d10v5_U73S5M
Xsky130_fd_pr__pfet_g5v0d10v5_PP2RNK_0 m1_790_6356# m1_779_5148# m1_n2158_9110# avdd
+ m1_790_6356# avdd m1_791_7588# m1_790_6356# m1_790_6356# m1_791_7588# avdd m1_790_6356#
+ m1_791_7588# m1_790_6356# m1_790_6356# m1_790_6356# m1_779_5148# m1_790_6356# m1_791_7588#
+ m1_791_7588# m1_n2158_9110# avdd m1_790_6356# m1_779_5148# m1_790_6356# m1_790_6356#
+ m1_n2158_9110# m1_791_7588# m1_3549_9621# avdd m1_n2158_9110# m1_790_6356# m1_790_6356#
+ m1_790_6356# m1_n2158_9110# m1_790_6356# m1_n2158_9110# m1_790_6356# m1_791_7588#
+ m1_790_6356# m1_n2158_9110# m1_n2158_9110# m1_790_6356# m1_791_7588# m1_790_6356#
+ avdd m1_n2158_9110# m1_3549_9621# avdd avdd sky130_fd_pr__pfet_g5v0d10v5_PP2RNK
Xsky130_fd_pr__nfet_g5v0d10v5_79TVLH_0 li_9924_630# m1_180_3630# li_9924_630# vinn
+ vinp m1_180_3630# m1_180_3630# li_9924_630# vinn li_9924_630# vinp li_9924_630#
+ vinn vinn vinn avss vinp li_9924_630# vinp m1_806_3964# vinn avss vinp li_9924_630#
+ li_9924_630# vinn vinp vinp m1_180_3630# m1_180_3630# li_9924_630# vinn vinn li_9924_630#
+ m1_806_3964# li_9924_630# vinn vinp m1_806_3964# m1_806_3964# avss vinp m1_180_3630#
+ vinp li_9924_630# vinp vinn m1_806_3964# m1_806_3964# vinp avss avss li_9924_630#
+ vinn sky130_fd_pr__nfet_g5v0d10v5_79TVLH
Xsky130_fd_pr__nfet_g5v0d10v5_2B7385_0 avss avss m1_n5910_1250# avss m1_n5910_1250#
+ m1_n5910_1250# m1_n5910_1250# m1_n5910_1250# avss avss m1_n5910_1250# avss avss
+ avss m1_n5910_1250# avss li_9924_630# li_9924_630# m1_n5910_1250# m1_n5910_1250#
+ m1_n5910_1250# li_9924_630# m1_n5910_1250# m1_n5910_1250# m1_n5910_1250# avss li_9924_630#
+ li_9924_630# avss m1_n5910_1250# m1_n5910_1250# avss m1_n5910_1250# avss li_9924_630#
+ li_9924_630# m1_n5910_1250# m1_n5910_1250# sky130_fd_pr__nfet_g5v0d10v5_2B7385
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_11 m1_n5904_n2678# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_79TVLH_1 li_9924_630# m1_806_3964# li_9924_630# vinp
+ vinn m1_806_3964# m1_806_3964# li_9924_630# vinp li_9924_630# vinn li_9924_630#
+ vinp vinp vinp avss vinn li_9924_630# vinn m1_180_3630# vinp avss vinn li_9924_630#
+ li_9924_630# vinp vinn vinn m1_806_3964# m1_806_3964# li_9924_630# vinp vinp li_9924_630#
+ m1_180_3630# li_9924_630# vinp vinn m1_180_3630# m1_180_3630# avss vinn m1_806_3964#
+ vinn li_9924_630# vinn vinp m1_180_3630# m1_180_3630# vinn avss avss li_9924_630#
+ vinp sky130_fd_pr__nfet_g5v0d10v5_79TVLH
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_12 m1_n5902_n1890# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_5X2ZTR_0 m1_790_6356# m1_n5902_n1100# m1_n5902_n1100#
+ m1_n5902_n1100# avss m1_n5906_n318# avss m1_n3947_7845# m1_23556_n2064# m1_n5902_n1100#
+ avss m1_n5902_n1100# avss m1_n5906_n318# m1_n5902_n1100# m1_n3947_7845# avss m1_n5902_n1100#
+ avss m1_22524_n1868# m1_n5906_n318# m1_23556_n2064# avss m1_n5902_n1100# m1_n3947_7845#
+ m1_n3947_7845# m1_n5902_n1100# m1_n5902_n1100# m1_22524_n1868# m1_n5906_n318# m1_790_6356#
+ m1_n5902_n1100# m1_n5902_n1100# avss m1_23556_n2064# m1_n5906_n318# m1_n5902_n1100#
+ m1_790_6356# m1_n5912_464# m1_n5902_n1100# m1_n5902_n1100# avss m1_22524_n1868#
+ avss m1_n5902_n1100# m1_180_4838# m1_23556_n2064# avss avss m1_22524_n1868# m1_n5902_n1100#
+ m1_n5902_n1100# m1_n5902_n1100# m1_790_6356# m1_n5902_n1100# m1_180_4838# avss avss
+ m1_n5902_n1100# m1_n5902_n1100# m1_22524_n1868# m1_23556_n2064# m1_n5902_n1100#
+ m1_n5902_n1100# m1_n5902_n1100# m1_180_4838# m1_180_4838# m1_n5902_n1100# m1_22524_n1868#
+ m1_n5902_n1100# m1_n5902_n1100# m1_n5902_n1100# m1_23556_n2064# m1_790_6356# m1_n5902_n1100#
+ m1_n5902_n1100# m1_n5902_n1100# m1_n5902_n1100# m1_n5906_n318# m1_n5902_n1100# m1_n3947_7845#
+ m1_180_4838# sky130_fd_pr__nfet_g5v0d10v5_5X2ZTR
Xsky130_fd_pr__nfet_g5v0d10v5_WK95DB_0 avss m1_n3080_8896# vb3 vb3 vb3 li_9924_630#
+ li_9924_630# vb3 vb3 m1_n3080_8896# m1_n3080_8896# vb3 vb3 li_9924_630# vb3 avss
+ m1_n3080_8896# avss avss avss m1_n3080_8896# li_9924_630# sky130_fd_pr__nfet_g5v0d10v5_WK95DB
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_13 m1_n5902_n1100# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14/a_50_n200#
+ avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_15 m1_n5910_1250# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_3QL9S5_0 m1_12142_11768# m1_n3334_8532# avdd m1_n3561_8311#
+ sky130_fd_pr__pfet_g5v0d10v5_3QL9S5
Xsky130_fd_pr__nfet_g5v0d10v5_PGZBW9_0 m1_n4694_n312# m1_n4694_n312# m1_n5902_n1890#
+ m1_n5902_n1890# avss m1_n4694_n312# avss m1_n4694_n312# m1_n4694_n312# avss m1_n4694_n312#
+ m1_n4694_n312# m1_n4694_n312# avss avss m1_n4694_n312# m1_n5904_n2678# m1_n4694_n312#
+ avss m1_n4694_n312# avss avss m1_n4694_n312# m1_n4694_n312# m1_n5902_n1890# avss
+ m1_n4694_n312# m1_n5902_n1890# m1_n4694_n312# m1_n4694_n312# m1_n5904_n2678# avss
+ avss m1_n4694_n312# m1_n4694_n312# m1_n5904_n2678# avss m1_n5904_n2678# m1_n4694_n312#
+ m1_n5902_n1890# avss m1_n4694_n312# m1_n4694_n312# m1_n4694_n312# m1_n5904_n2678#
+ m1_n4694_n312# m1_n5904_n2678# avss avss avss avss m1_n5902_n1890# avss m1_n4694_n312#
+ sky130_fd_pr__nfet_g5v0d10v5_PGZBW9
Xsky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD_1 avdd m1_n3264_4838# avdd m1_n3264_4838# avdd
+ m1_n3264_4838# avdd avdd avdd m1_n3264_4838# m1_n3667_4379# avdd avdd avdd m1_n3667_4379#
+ m1_n3667_4379# m1_n3667_4379# m1_n3667_4379# m1_n3667_4379# m1_n3264_4838# avdd
+ m1_n3264_4838# sky130_fd_pr__pfet_g5v0d10v5_U4Z9ZD
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_16 m1_n5912_464# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__res_generic_po_U7N8A7_0 avss avss m1_32006_n358# m1_32128_n282# m1_32714_1904#
+ m1_32128_n282# m1_32006_n358# m1_32250_1542# m1_32372_1542# vout avss m1_32250_1542#
+ avss m1_32494_n358# m1_32854_1648# m1_32616_n282# m1_32372_1542# m1_32616_n282#
+ vout avss m1_32494_n358# sky130_fd_pr__res_generic_po_U7N8A7
Xsky130_fd_pr__pfet_g5v0d10v5_3QL9S5_1 m1_12142_11768# m1_13086_11886# avdd m1_n3208_8640#
+ sky130_fd_pr__pfet_g5v0d10v5_3QL9S5
Xsky130_fd_pr__pfet_g5v0d10v5_QSKB8C_0 m1_n3947_7845# m1_n3947_7845# avdd m1_2256_n728#
+ m1_n3947_7845# m1_n3777_8065# m1_n3947_7845# m1_n4692_n1074# m1_n4692_n1074# m1_n3947_7845#
+ m1_n3947_7845# m1_n4182_7627# m1_25484_9858# m1_2256_n728# m1_n3947_7845# avdd m1_n3947_7845#
+ m1_n4704_472# m1_25484_9858# m1_n3947_7845# m1_n3947_7845# m1_n4692_n1074# m1_n3947_7845#
+ m1_n3947_7845# m1_n4182_7627# m1_n3947_7845# m1_n3947_7845# avdd m1_25484_9858#
+ avdd avdd m1_n3947_7845# m1_25484_9858# m1_23420_9858# m1_n3947_7845# m1_n3947_7845#
+ m1_n4692_n1074# m1_n3947_7845# m1_n3947_7845# avdd avdd m1_n3947_7845# avdd m1_23420_9858#
+ avdd m1_n4704_472# m1_n3947_7845# m1_n3947_7845# avdd m1_n3947_7845# m1_n4182_7627#
+ m1_n4692_n1074# avdd m1_n3947_7845# m1_n3947_7845# m1_n3947_7845# avdd m1_25484_9858#
+ m1_n3947_7845# m1_n3947_7845# m1_25484_9858# m1_n4692_n1074# m1_2256_n728# avdd
+ m1_n4704_472# avdd m1_n3947_7845# m1_n3777_8065# m1_n3947_7845# m1_n3777_8065# m1_n4692_n1074#
+ m1_23420_9858# m1_n3947_7845# m1_n3947_7845# m1_n3947_7845# m1_n4704_472# m1_2256_n728#
+ m1_n3947_7845# sky130_fd_pr__pfet_g5v0d10v5_QSKB8C
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_17 m1_n5906_n318# avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__pfet_g5v0d10v5_QRKB8C_0 m1_n3777_8065# m1_n3777_8065# avdd m1_23420_9858#
+ m1_n3777_8065# avdd avdd m1_n3777_8065# m1_n3777_8065# avdd m1_n3777_8065# avdd
+ avdd m1_n4182_7627# m1_n3777_8065# m1_n3777_8065# avdd m1_25484_9858# avdd avdd
+ avdd m1_25484_9858# m1_n3777_8065# avdd avdd m1_n3777_8065# m1_n3777_8065# avdd
+ m1_n3777_8065# m1_n3777_8065# m1_23420_9858# avdd avdd avdd m1_23420_9858# m1_25484_9858#
+ m1_n3777_8065# m1_n3777_8065# avdd m1_n3777_8065# avdd avdd m1_n3777_8065# m1_n4182_7627#
+ m1_n3777_8065# m1_n3777_8065# m1_n4182_7627# avdd m1_n4182_7627# m1_n3777_8065#
+ m1_n3777_8065# m1_n3777_8065# m1_n3777_8065# avdd m1_n3777_8065# m1_n3777_8065#
+ avdd m1_25484_9858# avdd m1_n3777_8065# m1_25484_9858# m1_n3777_8065# m1_n3777_8065#
+ avdd m1_n3777_8065# avdd m1_n3777_8065# avdd avdd m1_n3777_8065# m1_n3777_8065#
+ m1_25484_9858# m1_23420_9858# m1_n3777_8065# sky130_fd_pr__pfet_g5v0d10v5_QRKB8C
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18/a_50_n200#
+ avss avss m1_n6000_2704# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__cap_mim_m3_1_Z5XS7R_1 m1_16202_3432# m1_n592_3104# m1_32854_1648# m1_16202_3432#
+ m1_32714_1904# m1_32714_1904# m1_n592_3104# m1_16202_3432# m1_32714_1904# m1_32854_1648#
+ m1_32854_1648# m1_n592_3104# sky130_fd_pr__cap_mim_m3_1_Z5XS7R
Xsky130_fd_pr__pfet_g5v0d10v5_EVM3FM_0 m1_790_6356# m1_790_6356# m1_790_6356# m1_n5910_1250#
+ m1_790_6356# m1_790_6356# m1_n2158_9110# m1_790_6356# avdd m1_790_6356# m1_n2158_9110#
+ m1_790_6356# avdd m1_n5910_1250# avdd avdd m1_n2158_9110# m1_n5910_1250# m1_n5910_1250#
+ avdd m1_n2158_9110# m1_n2158_9110# sky130_fd_pr__pfet_g5v0d10v5_EVM3FM
Xsky130_fd_pr__nfet_g5v0d10v5_CTEUHA_19 avss avss m1_n6000_2704# m1_n3667_4379# sky130_fd_pr__nfet_g5v0d10v5_CTEUHA
Xsky130_fd_pr__nfet_g5v0d10v5_DL2ZHN_0 m1_n5906_n318# m1_n5912_464# m1_n5912_464#
+ m1_n5912_464# avss m1_n5912_464# m1_23556_n2064# avss avss m1_n5912_464# m1_n5912_464#
+ avss m1_n5912_464# m1_22524_n1868# m1_n5906_n318# m1_n5912_464# m1_n5912_464# avss
+ avss avss m1_n5912_464# m1_n5912_464# m1_n5906_n318# m1_23556_n2064# m1_n5912_464#
+ m1_n5912_464# avss avss m1_n5906_n318# m1_n5912_464# m1_n5912_464# avss avss m1_n5912_464#
+ m1_22524_n1868# m1_22524_n1868# m1_n5912_464# m1_n5912_464# avss m1_n5906_n318#
+ m1_n5912_464# m1_23556_n2064# avss m1_n5912_464# avss avss m1_n5912_464# m1_n5912_464#
+ m1_23556_n2064# m1_n5912_464# m1_n5906_n318# m1_n5912_464# m1_22524_n1868# avss
+ m1_n5912_464# avss avss avss m1_n5912_464# m1_n5912_464# m1_23556_n2064# m1_n5912_464#
+ avss avss m1_n5912_464# m1_n5912_464# avss avss m1_23556_n2064# avss m1_n5912_464#
+ m1_n5912_464# m1_n5912_464# avss avss m1_22524_n1868# m1_22524_n1868# avss sky130_fd_pr__nfet_g5v0d10v5_DL2ZHN
Xsky130_fd_pr__pfet_g5v0d10v5_Q46EE6_0 m1_n3445_8429# m1_n3334_8532# m1_n3334_8532#
+ avdd m1_n3561_8311# m1_n3334_8532# m1_n3445_8429# m1_n3208_8640# avdd m1_n3445_8429#
+ avdd avdd m1_n3334_8532# m1_n3445_8429# avdd m1_n3208_8640# m1_n3334_8532# m1_n5902_n1100#
+ m1_n5902_n1100# m1_n3334_8532# avdd m1_n3334_8532# m1_n5902_n1100# m1_n5902_n1100#
+ m1_n3334_8532# avdd m1_n3334_8532# avdd m1_n5902_n1100# m1_n3334_8532# sky130_fd_pr__pfet_g5v0d10v5_Q46EE6
Xsky130_fd_pr__nfet_g5v0d10v5_UGZTXE_0 vb3 vb3 m1_n4694_n312# m1_16202_3432# m1_n5902_n1890#
+ avss vb3 m1_n5904_n2678# vb3 vb3 m1_n5902_n1890# vb3 vb3 vb3 avss m1_n5904_n2678#
+ avss vb3 m1_n4694_n312# vb3 m1_16202_3432# vb3 avss m1_n5904_n2678# vb3 vb3 m1_16202_3432#
+ m1_n5902_n1890# avss m1_n4694_n312# vb3 vb3 m1_n4694_n312# m1_n5904_n2678# m1_n5902_n1890#
+ vb3 vb3 avss m1_16202_3432# vb3 avss m1_n4694_n312# vb3 m1_n4694_n312# m1_n5902_n1890#
+ avss vb3 vb3 m1_16202_3432# vb3 m1_16202_3432# m1_n4694_n312# vb3 m1_n5904_n2678#
+ m1_n5904_n2678# m1_16202_3432# m1_n5902_n1890# vb3 sky130_fd_pr__nfet_g5v0d10v5_UGZTXE
Xsky130_fd_pr__pfet_g5v0d10v5_XW23Q2_0 m1_779_5148# m1_791_7588# m1_3549_9621# m1_779_5148#
+ avdd avdd m1_779_5148# m1_779_5148# avdd m1_779_5148# avdd m1_779_5148# m1_779_5148#
+ m1_779_5148# avdd m1_779_5148# avdd avdd m1_791_7588# m1_779_5148# m1_791_7588#
+ m1_779_5148# m1_779_5148# m1_791_7588# avdd avdd m1_779_5148# m1_791_7588# m1_779_5148#
+ m1_779_5148# avdd m1_791_7588# m1_779_5148# m1_3549_9621# m1_779_5148# avdd m1_779_5148#
+ avdd m1_791_7588# avdd avdd m1_779_5148# avdd m1_791_7588# avdd m1_779_5148# sky130_fd_pr__pfet_g5v0d10v5_XW23Q2
Xsky130_fd_pr__nfet_g5v0d10v5_HG2LSW_0 vb3 vb3 avss avss sky130_fd_pr__nfet_g5v0d10v5_HG2LSW
Xsky130_fd_pr__nfet_g5v0d10v5_N64HU4_0 avss avss avss avss ibias m1_n3955_n943# m1_n3955_n943#
+ avss m1_n4700_n2510# m1_n4700_n2510# m1_n4700_n2510# m1_n4685_n1863# m1_n3955_n943#
+ m1_n3955_n943# m1_n3955_n943# m1_n3955_n943# m1_n3561_8311# m1_n3955_n943# m1_n3955_n943#
+ m1_282_n2232# m1_n3955_n943# m1_n3561_8311# m1_n3955_n943# m1_n3561_8311# m1_n4700_n2510#
+ m1_n3561_8311# avss avss avss m1_n3561_8311# m1_n3955_n943# m1_n3955_n943# m1_n4685_n1863#
+ m1_n4700_n2510# sky130_fd_pr__nfet_g5v0d10v5_N64HU4
Xsky130_fd_pr__nfet_g5v0d10v5_RMXH5H_0 m1_18790_1436# avss m1_n4704_472# m1_n4704_472#
+ avss m1_18790_1436# m1_18790_1436# m1_n4704_472# avss avss avss m1_18790_1436# avss
+ avss avss m1_n4704_472# m1_18790_1436# m1_n4704_472# m1_18790_1436# m1_18790_1436#
+ m1_18790_1436# avss avss m1_n4704_472# m1_n4704_472# avss sky130_fd_pr__nfet_g5v0d10v5_RMXH5H
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_10 m1_n3208_8640# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_TT9EEV_0 m1_n1154_3624# avdd avdd m1_16202_3432# m1_180_4838#
+ m1_180_4838# m1_n1154_3624# m1_180_4838# m1_n4694_n312# avdd m1_n1154_3624# m1_16202_3432#
+ avdd avdd m1_180_4838# avdd m1_180_4838# m1_n1154_3624# m1_n4694_n312# m1_n592_3104#
+ m1_180_4838# m1_180_4838# avdd m1_n4694_n312# m1_180_4838# m1_n592_3104# avdd m1_180_4838#
+ sky130_fd_pr__pfet_g5v0d10v5_TT9EEV
Xsky130_fd_pr__pfet_g5v0d10v5_BH2H9S_0 m1_n3080_8896# m1_n3080_8896# m1_n2158_9110#
+ avdd m1_n3080_8896# avdd m1_n3080_8896# m1_n2158_9110# m1_n3080_8896# m1_n3080_8896#
+ avdd m1_n2158_9110# m1_n3080_8896# avdd avdd m1_n3080_8896# m1_n3080_8896# m1_n3080_8896#
+ m1_n3080_8896# avdd m1_n2158_9110# avdd m1_n3080_8896# m1_n3080_8896# m1_n3080_8896#
+ m1_n3080_8896# avdd avdd avdd avdd m1_n3080_8896# avdd avdd m1_n2158_9110# avdd
+ m1_n3080_8896# m1_n3080_8896# m1_n2158_9110# sky130_fd_pr__pfet_g5v0d10v5_BH2H9S
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_11 m1_n3334_8532# avdd m1_n1846_3922# avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__nfet_g5v0d10v5_NMXZ6U_0 m1_n4700_n2510# m1_n4698_n3450# avss m1_n4700_n2510#
+ m1_n4698_n3450# m1_n4698_n3450# avss avss avss avss m1_n4698_n3450# avss m1_n4698_n3450#
+ m1_n4698_n3450# m1_n4700_n2510# m1_n4698_n3450# m1_n4698_n3450# avss m1_n4698_n3450#
+ m1_n4700_n2510# m1_n4698_n3450# m1_n4700_n2510# avss m1_n4685_n1863# m1_n4698_n3450#
+ m1_n4700_n2510# m1_n4698_n3450# avss avss avss sky130_fd_pr__nfet_g5v0d10v5_NMXZ6U
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_12 avdd avdd m1_n1846_3922# m1_n3947_7845# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_14 avdd avdd m1_n1846_3922# m1_n3445_8429# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
Xsky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13 avdd avdd m1_n1846_3922# m1_n592_3104# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD
C0 m1_n1846_3922# m1_779_5148# 0.523504f
C1 m1_n6000_2704# m1_n5902_n1100# 0.210379f
C2 m1_779_5148# m1_n2158_9110# 0.881995f
C3 m1_n4694_n312# m1_n4704_472# 1.908395f
C4 m1_n3667_4379# m1_n3264_4838# 3.886719f
C5 m1_n1154_3624# m1_n592_3104# 0.554139f
C6 m1_n4694_n312# m1_n4698_n3450# 0.162463f
C7 m1_n5910_1250# m1_n4704_472# 1.887962f
C8 m1_790_6356# m1_n592_3104# 19.510752f
C9 m1_n1154_3624# m1_n4692_n1074# 0.236899f
C10 m1_n9267_3854# avdd 0.105765f
C11 m1_n3080_8896# m1_n4692_n1074# 0.185369f
C12 m1_n5904_n2678# m1_n5902_n1100# 1.8423f
C13 m1_n3264_4838# m1_n4704_472# 0.11444f
C14 m1_13086_11886# m1_n3208_8640# 0.511976f
C15 m1_n6000_2704# m1_n4685_n1863# 0.179503f
C16 m1_790_6356# m1_16202_3432# 0.273673f
C17 m1_790_6356# m1_n4692_n1074# 1.88212f
C18 m1_n3334_8532# m1_790_6356# 1.865219f
C19 m1_180_4838# m1_n592_3104# 3.81405f
C20 m1_n1154_3624# m1_180_3630# 24.285135f
C21 m1_n3080_8896# m1_180_3630# 0.130359f
C22 m1_180_4838# m1_16202_3432# 3.612051f
C23 m1_180_3630# m1_790_6356# 23.124596f
C24 m1_n4700_n2510# m1_n4694_n312# 0.260656f
C25 m1_n1154_3624# m1_n4704_472# 2.902205f
C26 m1_23556_n2064# m1_n5906_n318# 3.373696f
C27 m1_n3561_8311# m1_791_7588# 0.510596f
C28 m1_2256_n728# m1_n2158_9110# 0.164043f
C29 vb3 net12 10.246552f
C30 m1_790_6356# m1_n4704_472# 0.82824f
C31 m1_180_4838# m1_180_3630# 0.715597f
C32 vinn m1_n592_3104# 5.82961f
C33 vout m1_n5902_n1100# 0.76128f
C34 m1_3549_9621# m1_779_5148# 2.131759f
C35 ibias vinn 0.943112f
C36 m1_n6000_2704# m1_n9267_3854# 0.197128f
C37 m1_180_4838# m1_n4704_472# 1.242579f
C38 m1_32854_1648# avdd 0.394939f
C39 m1_n8442_3847# dvdd 0.103652f
C40 net12 net29 2.181938f
C41 avdd m1_n592_3104# 0.124089p
C42 m1_n3667_4379# vinn 0.110177f
C43 m1_n5902_n1890# m1_n5902_n1100# 0.809929f
C44 ibias avdd 0.686189f
C45 m1_n3561_8311# m1_n3208_8640# 2.824089f
C46 vb3 net29 2.171696f
C47 m1_18668_3467# m1_180_4838# 1.381749f
C48 m1_13086_11886# m1_790_6356# 0.353704f
C49 vinn m1_180_3630# 0.668658f
C50 avdd m1_n4692_n1074# 11.476912f
C51 avdd m1_16202_3432# 1.242312f
C52 avdd m1_n3334_8532# 9.987501f
C53 m1_n3667_4379# avdd 3.479839f
C54 m1_n1154_3624# m1_806_3964# 13.923638f
C55 net12 li_9924_630# -2.243941f
C56 m1_n3947_7845# vinp 0.145761f
C57 vinn m1_n4704_472# 0.381894f
C58 avdd m1_180_3630# 15.279448f
C59 m1_806_3964# m1_790_6356# 20.376215f
C60 m1_n3561_8311# m1_n5910_1250# 1.120438f
C61 vb3 li_9924_630# 13.9456f
C62 m1_18790_1436# m1_16202_3432# 0.177436f
C63 m1_23420_9858# m1_n3947_7845# 2.928139f
C64 avdd m1_n4704_472# 10.358822f
C65 m1_180_4838# m1_806_3964# 0.204417f
C66 m1_2256_n728# m1_3549_9621# 0.101797f
C67 m1_18668_3467# avdd 4.027752f
C68 m1_n4182_7627# m1_n4704_472# -0.748629f
C69 ibias m1_n6000_2704# 0.150379f
C70 m1_n9267_3854# ena 0.105639f
C71 m1_n3561_8311# m1_n1154_3624# 0.852564f
C72 m1_n6000_2704# m1_n4692_n1074# 0.175739f
C73 m1_n3561_8311# m1_n3080_8896# 1.985486f
C74 m1_18790_1436# m1_n4704_472# 0.855844f
C75 m1_n3667_4379# m1_n6000_2704# 0.932488f
C76 m1_n3561_8311# m1_790_6356# 2.316047f
C77 m1_13086_11886# avdd 5.568506f
C78 vinn m1_806_3964# 10.835169f
C79 m1_2256_n728# m1_779_5148# 0.126477f
C80 m1_32714_1904# m1_n3947_7845# 0.227724f
C81 vb3 m1_n8442_3847# 0.242026f
C82 m1_n1846_3922# m1_n592_3104# 1.049568f
C83 avdd m1_806_3964# 6.125107f
C84 m1_n5904_n2678# m1_16202_3432# -2.333696f
C85 m1_n6000_2704# m1_n4704_472# 0.185922f
C86 m1_n3561_8311# m1_n3777_8065# 6.719668f
C87 m1_n1846_3922# m1_n3334_8532# 0.464791f
C88 m1_n4692_n1074# m1_n2158_9110# 0.354185f
C89 m1_n6000_2704# m1_n4698_n3450# 0.183464f
C90 m1_180_3630# m1_n5904_n2678# 1.74053f
C91 m1_n1846_3922# m1_180_3630# 0.712613f
C92 m1_180_3630# m1_n2158_9110# 2.57189f
C93 m1_n5904_n2678# m1_n4704_472# 0.582905f
C94 net12 net28 0.758131f
C95 li_9924_630# vinp 11.733767f
C96 vout m1_n592_3104# 67.67779f
C97 m1_790_6356# m1_23556_n2064# -0.552379f
C98 vb3 net28 2.169403f
C99 m1_n3561_8311# avdd 21.248497f
C100 m1_n6000_2704# m1_n4700_n2510# 0.212934f
C101 vout m1_16202_3432# 29.575033f
C102 m1_n6000_2704# m1_n5912_464# 0.474654f
C103 vb3 m1_n4694_n312# 7.651504f
C104 m1_12142_11768# m1_n3334_8532# 0.615444f
C105 vb3 m1_n5910_1250# 0.388623f
C106 vout m1_n4704_472# 0.489022f
C107 m1_n3947_7845# m1_n3777_8065# 14.542556f
C108 m1_n5902_n1890# m1_180_3630# 0.585099f
C109 m1_806_3964# m1_n5904_n2678# 6.430725f
C110 m1_n3445_8429# m1_n3208_8640# 1.994293f
C111 m1_3549_9621# m1_n4692_n1074# 0.452149f
C112 m1_n1846_3922# m1_806_3964# 0.512479f
C113 m1_25484_9858# m1_n3777_8065# 6.079924f
C114 m1_806_3964# m1_n2158_9110# 0.417818f
C115 m1_n5902_n1890# m1_n4704_472# 0.445875f
C116 vout m1_22524_n1868# 0.292619f
C117 vb3 m1_n1154_3624# 0.401852f
C118 vb3 m1_n3080_8896# 4.932774f
C119 li_9924_630# m1_n5910_1250# 8.92591f
C120 m1_779_5148# m1_n4692_n1074# 4.09055f
C121 avdd m1_n3947_7845# 17.378897f
C122 vout m1_n5912_464# 0.958703f
C123 m1_12142_11768# m1_13086_11886# 0.397736f
C124 m1_n3561_8311# m1_n1846_3922# 0.479564f
C125 m1_25484_9858# avdd 1.28985f
C126 m1_n3561_8311# m1_n2158_9110# 0.130372f
C127 m1_180_3630# m1_779_5148# 0.723394f
C128 m1_n4182_7627# m1_n3947_7845# 13.333585f
C129 m1_n5902_n1890# m1_806_3964# 0.492921f
C130 m1_n5902_n1100# m1_n592_3104# 0.112606f
C131 m1_282_n2232# m1_n3955_n943# 0.268666f
C132 m1_25484_9858# m1_n4182_7627# 1.892255f
C133 li_9924_630# m1_n3080_8896# -1.940126f
C134 m1_n5902_n1100# m1_16202_3432# 0.31357f
C135 m1_n3334_8532# m1_n5902_n1100# 2.49195f
C136 vb3 vinn 0.613709f
C137 m1_n3955_n943# m1_2256_n728# 0.595747f
C138 m1_2256_n728# m1_n592_3104# 0.130321f
C139 m1_n3445_8429# m1_n3777_8065# 0.172941f
C140 m1_180_3630# m1_n5902_n1100# 0.426331f
C141 m1_n3955_n943# m1_n4685_n1863# 0.392301f
C142 m1_2256_n728# m1_n4692_n1074# 10.169897f
C143 m1_n8442_3847# m1_n3264_4838# 0.52173f
C144 m1_180_4838# m1_n5906_n318# -0.555734f
C145 m1_n5902_n1100# m1_n4704_472# 0.103718f
C146 m1_n5910_1250# m1_791_7588# 0.248648f
C147 m1_n4685_n1863# m1_n4692_n1074# 0.122713f
C148 m1_n3561_8311# m1_12142_11768# 1.037745f
C149 m1_2256_n728# m1_180_3630# 0.509775f
C150 m1_n1154_3624# vinp 0.572779f
C151 m1_806_3964# m1_779_5148# 0.366362f
C152 dvdd ena 0.540205f
C153 net28 m1_n4694_n312# 0.582207f
C154 m1_n1846_3922# m1_n3947_7845# 0.59511f
C155 li_9924_630# vinn 11.322492f
C156 m1_2256_n728# m1_n4704_472# 0.220238f
C157 m1_n5902_n1100# m1_22524_n1868# 3.858514f
C158 avdd m1_n3445_8429# 8.188938f
C159 m1_n4685_n1863# m1_n3750_n668# 0.360933f
C160 m1_n6000_2704# net12 0.203506f
C161 m1_n3080_8896# m1_791_7588# 0.13079f
C162 m1_180_4838# vinp 4.534452f
C163 m1_n5910_1250# m1_n3208_8640# 2.4961f
C164 vb3 m1_n6000_2704# 0.554873f
C165 ibias m1_n9267_3854# 0.181597f
C166 m1_790_6356# m1_791_7588# 14.444685f
C167 m1_n4685_n1863# m1_n4698_n3450# 2.519198f
C168 m1_n5912_464# m1_n5902_n1100# 0.565285f
C169 m1_282_n2232# m1_n4700_n2510# 0.105474f
C170 m1_n3667_4379# m1_n9267_3854# 0.526141f
C171 m1_n3561_8311# m1_779_5148# 1.420192f
C172 net12 m1_n5904_n2678# 5.639711f
C173 m1_23420_9858# m1_n3777_8065# 4.126304f
C174 m1_n5910_1250# m1_n3264_4838# 0.217356f
C175 vb3 m1_n5904_n2678# 8.226118f
C176 vinn vinp 9.772527f
C177 m1_n3080_8896# m1_n3208_8640# 1.519337f
C178 m1_2256_n728# m1_806_3964# 1.524994f
C179 m1_n1154_3624# m1_n4694_n312# -0.843515f
C180 m1_n8442_3847# vinn 0.192501f
C181 vb3 m1_n1846_3922# 0.244264f
C182 m1_n9267_3854# m1_n4704_472# 0.150144f
C183 m1_n3208_8640# m1_790_6356# 0.46204f
C184 m1_n4685_n1863# m1_n4700_n2510# 0.982989f
C185 avdd vinp 11.533832f
C186 m1_32854_1648# m1_n592_3104# 0.586444f
C187 m1_n8442_3847# avdd 0.173938f
C188 m1_n5910_1250# m1_n3080_8896# 5.603479f
C189 m1_n6000_2704# m1_n5906_n318# 0.206979f
C190 m1_180_4838# m1_n4694_n312# 2.597208f
C191 m1_n4182_7627# vinp 0.164168f
C192 m1_23420_9858# avdd 2.60346f
C193 ibias m1_n3955_n943# 1.169057f
C194 m1_32854_1648# m1_16202_3432# 0.6408f
C195 m1_n5910_1250# m1_790_6356# 7.976317f
C196 avdd m1_791_7588# 1.210982f
C197 m1_n592_3104# m1_n4692_n1074# 0.137222f
C198 m1_16202_3432# m1_n592_3104# 5.813296f
C199 m1_n1846_3922# m1_n3445_8429# 0.420794f
C200 ibias m1_n4692_n1074# 0.212011f
C201 m1_23420_9858# m1_n4182_7627# 3.388911f
C202 m1_n3561_8311# m1_2256_n728# 2.97024f
C203 ibias m1_n3667_4379# 0.154113f
C204 m1_180_3630# m1_n592_3104# -3.151957f
C205 vb3 m1_n5902_n1890# 7.836075f
C206 m1_n1154_3624# m1_790_6356# 21.520802f
C207 m1_n3955_n943# m1_n3750_n668# 0.340553f
C208 m1_180_3630# m1_n4692_n1074# 1.994658f
C209 m1_n3080_8896# m1_790_6356# 0.105232f
C210 m1_n592_3104# m1_n4704_472# 6.296457f
C211 ibias m1_n3750_n668# 0.437225f
C212 avdd m1_n3208_8640# 7.662561f
C213 m1_n6000_2704# m1_n8442_3847# 0.361847f
C214 m1_32714_1904# avdd 1.923648f
C215 m1_n3955_n943# m1_n4698_n3450# 0.264084f
C216 avdd m1_n4694_n312# 0.765742f
C217 m1_n1154_3624# m1_180_4838# 9.55744f
C218 m1_n4692_n1074# m1_n4704_472# 2.01833f
C219 m1_16202_3432# m1_n4704_472# 1.594152f
C220 m1_n5902_n1100# m1_23556_n2064# 2.778417f
C221 m1_18668_3467# m1_n592_3104# 0.184357f
C222 m1_n4698_n3450# m1_n4692_n1074# 1.913527f
C223 m1_180_4838# m1_790_6356# 2.541534f
C224 m1_n5904_n2678# vinp 19.253344f
C225 m1_180_3630# m1_n4704_472# 1.92039f
C226 m1_n5910_1250# avdd 10.953123f
C227 m1_n3947_7845# m1_n5902_n1100# 3.591318f
C228 m1_n1846_3922# vinp 0.273767f
C229 vout m1_n5906_n318# 0.251261f
C230 avdd m1_n3264_4838# 2.927261f
C231 vinp m1_n2158_9110# 21.00029f
C232 vinn m1_n1154_3624# 0.153798f
C233 m1_13086_11886# m1_n3334_8532# 1.576239f
C234 m1_n3955_n943# m1_n4700_n2510# 1.264596f
C235 m1_n3750_n668# m1_n4698_n3450# 0.312309f
C236 vb3 m1_779_5148# 2.38452f
C237 m1_2256_n728# m1_n3947_7845# 2.932078f
C238 m1_n1846_3922# m1_791_7588# 0.410755f
C239 m1_791_7588# m1_n2158_9110# -4.560299f
C240 m1_n4700_n2510# m1_n4692_n1074# 0.112312f
C241 avdd m1_n1154_3624# 72.935555f
C242 m1_13086_11886# m1_180_3630# 0.233319f
C243 m1_n6000_2704# m1_n4694_n312# 0.287221f
C244 m1_806_3964# m1_n4692_n1074# 0.578376f
C245 m1_n3080_8896# avdd 40.05257f
C246 vinn m1_180_4838# 0.606327f
C247 avdd m1_790_6356# 19.970827f
C248 net29 m1_779_5148# -0.571569f
C249 m1_n9267_3854# dvdd 0.608914f
C250 net12 m1_n5902_n1100# 4.90079f
C251 m1_180_3630# m1_806_3964# 5.347499f
C252 m1_n6000_2704# m1_n5910_1250# 0.835109f
C253 avdd m1_180_4838# 6.225294f
C254 m1_n5902_n1890# vinp 1.547996f
C255 m1_n4694_n312# m1_n5904_n2678# 7.503953f
C256 m1_n1846_3922# m1_n3208_8640# 0.400037f
C257 avdd m1_n3777_8065# 33.530792f
C258 m1_806_3964# m1_n4704_472# 1.99496f
C259 m1_n3561_8311# m1_n3955_n943# 5.296822f
C260 li_9924_630# m1_779_5148# 0.170767f
C261 m1_n4700_n2510# m1_n4698_n3450# 1.772426f
C262 m1_n3561_8311# m1_n4692_n1074# 0.113181f
C263 m1_n4182_7627# m1_n3777_8065# 3.521509f
C264 m1_n3561_8311# m1_n3334_8532# 0.454196f
C265 vb3 m1_2256_n728# 0.862216f
C266 m1_n5912_464# m1_22524_n1868# 2.457647f
C267 m1_n5910_1250# m1_n1846_3922# 0.123067f
C268 avdd vinn 4.797814f
C269 m1_n5910_1250# m1_n2158_9110# -3.404715f
C270 m1_n3561_8311# m1_180_3630# 0.438931f
C271 m1_n1846_3922# m1_n3264_4838# 0.878571f
C272 m1_n3445_8429# m1_n5902_n1100# -0.448167f
C273 m1_3549_9621# m1_791_7588# 1.174547f
C274 m1_n1154_3624# m1_n5904_n2678# 1.805144f
C275 m1_n5902_n1100# m1_n5906_n318# 12.324423f
C276 m1_n1846_3922# m1_n1154_3624# 0.591179f
C277 vinp m1_779_5148# 0.253037f
C278 avdd m1_n4182_7627# 17.088707f
C279 m1_n3080_8896# m1_n1846_3922# 0.406765f
C280 m1_12142_11768# m1_n3208_8640# 0.45921f
C281 m1_n3080_8896# m1_n2158_9110# 17.28071f
C282 m1_n4694_n312# m1_n5902_n1890# 10.217694f
C283 m1_2256_n728# li_9924_630# 0.510869f
C284 m1_n1846_3922# m1_790_6356# 0.52304f
C285 m1_790_6356# m1_n2158_9110# 22.029453f
C286 m1_32854_1648# m1_n3947_7845# 0.193204f
C287 vb3 m1_n9267_3854# 0.145737f
C288 m1_779_5148# m1_791_7588# 13.407484f
C289 m1_n6000_2704# vinn 0.107124f
C290 m1_n3947_7845# m1_n592_3104# 1.305463f
C291 m1_n1846_3922# m1_180_4838# 0.552461f
C292 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18/a_50_n200# m1_n6000_2704# 0.17739f
C293 m1_n1846_3922# m1_n3777_8065# 0.548189f
C294 m1_n3947_7845# m1_n4692_n1074# 6.516981f
C295 m1_n3561_8311# m1_n4700_n2510# -0.126873f
C296 m1_n3947_7845# m1_16202_3432# 0.778141f
C297 m1_n6000_2704# avdd 0.285385f
C298 m1_25484_9858# m1_n4692_n1074# -1.488901f
C299 vout m1_790_6356# 0.246282f
C300 vinn m1_n5904_n2678# 0.790447f
C301 m1_n1846_3922# vinn 0.252776f
C302 vinn m1_n2158_9110# 20.958448f
C303 m1_n3947_7845# m1_n4704_472# 3.401505f
C304 vout m1_180_4838# 0.332375f
C305 avdd m1_n5904_n2678# 6.948539f
C306 m1_22524_n1868# m1_23556_n2064# 0.749358f
C307 m1_12142_11768# m1_790_6356# 0.546464f
C308 m1_n1846_3922# avdd 10.241329f
C309 m1_2256_n728# m1_23420_9858# -0.753585f
C310 avdd m1_n2158_9110# 9.76134f
C311 m1_2256_n728# m1_791_7588# 0.505947f
C312 net12 m1_n4692_n1074# 7.619293f
C313 m1_n5910_1250# m1_779_5148# 2.416432f
C314 m1_180_4838# m1_n5902_n1890# 0.101783f
C315 m1_n3947_7845# m1_22524_n1868# -0.537066f
C316 m1_n1846_3922# m1_n4182_7627# 0.548188f
C317 m1_3549_9621# m1_790_6356# 3.349084f
C318 vb3 m1_n4692_n1074# 2.700586f
C319 vb3 m1_16202_3432# 6.984681f
C320 m1_n5912_464# m1_23556_n2064# 2.949108f
C321 m1_n3667_4379# vb3 0.274202f
C322 m1_n4694_n312# m1_n5902_n1100# 2.0776f
C323 vb3 m1_180_3630# 0.202157f
C324 net29 m1_n4692_n1074# 2.431832f
C325 vinn m1_n5902_n1890# 18.731585f
C326 avdd vout -19.690844f
C327 m1_n3080_8896# m1_779_5148# 0.41781f
C328 m1_n6000_2704# m1_n5904_n2678# 0.232469f
C329 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14/a_50_n200# m1_n6000_2704# 0.184804f
C330 vb3 m1_n4704_472# 0.871242f
C331 m1_n8442_3847# m1_n9267_3854# 0.847881f
C332 m1_790_6356# m1_779_5148# 3.83268f
C333 m1_n3955_n943# li_9924_630# 0.489393f
C334 m1_n3334_8532# m1_n3445_8429# 13.860621f
C335 avdd m1_n5902_n1890# 3.039456f
C336 m1_n4685_n1863# m1_n4694_n312# 0.108618f
C337 m1_12142_11768# avdd 1.066746f
C338 m1_180_4838# m1_779_5148# 0.10895f
C339 li_9924_630# m1_n4692_n1074# 0.413052f
C340 m1_3549_9621# avdd 0.368962f
C341 li_9924_630# m1_180_3630# 1.916226f
C342 m1_n5904_n2678# m1_n2158_9110# 2.452492f
C343 m1_n5902_n1100# m1_790_6356# 8.963762f
C344 vinn m1_779_5148# 0.540778f
C345 m1_2256_n728# m1_n1154_3624# 0.569803f
C346 m1_2256_n728# m1_n3080_8896# 0.161154f
C347 m1_180_4838# m1_n5902_n1100# 3.823886f
C348 vinp m1_n592_3104# 0.120644f
C349 ibias vinp 0.315497f
C350 m1_n6000_2704# m1_n5902_n1890# 0.230754f
C351 m1_2256_n728# m1_790_6356# 1.731076f
C352 avdd m1_779_5148# 34.3809f
C353 ibias m1_n8442_3847# 0.153071f
C354 m1_13086_11886# m1_n3445_8429# 1.754364f
C355 m1_n5910_1250# m1_n9267_3854# 0.436556f
C356 m1_22524_n1868# m1_n5906_n318# 3.712793f
C357 m1_n3667_4379# m1_n8442_3847# 0.34374f
C358 m1_180_3630# vinp 11.012436f
C359 m1_n9267_3854# m1_n3264_4838# 0.159282f
C360 m1_791_7588# m1_n4692_n1074# 0.653221f
C361 m1_n5902_n1890# m1_n5904_n2678# 13.695122f
C362 m1_n3334_8532# m1_791_7588# 0.158251f
C363 vinp m1_n4704_472# 0.146426f
C364 li_9924_630# m1_806_3964# 3.424842f
C365 m1_n5902_n1890# m1_n2158_9110# 4.251904f
C366 avdd m1_n5902_n1100# 8.107554f
C367 m1_n5912_464# m1_n5906_n318# 14.035233f
C368 m1_32714_1904# m1_32854_1648# 7.996289f
C369 m1_32714_1904# m1_n592_3104# 0.556922f
C370 net28 m1_n4692_n1074# 3.781344f
C371 ibias m1_n4694_n312# 0.165171f
C372 m1_2256_n728# avdd 9.947802f
C373 m1_n3334_8532# m1_n3208_8640# 12.10555f
C374 m1_25484_9858# m1_n3947_7845# 5.1524f
C375 m1_32714_1904# m1_16202_3432# 5.23945f
C376 m1_n3561_8311# m1_n3445_8429# 11.666098f
C377 m1_n4694_n312# m1_n4692_n1074# 6.608271f
C378 m1_n4694_n312# m1_16202_3432# 2.223908f
C379 m1_n3955_n943# m1_n5910_1250# 0.15611f
C380 m1_n3561_8311# li_9924_630# 0.113562f
C381 ibias m1_n5910_1250# 0.125541f
C382 m1_806_3964# vinp 1.175008f
C383 m1_n3445_8429# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.648804f
C384 m1_n4700_n2510# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 6.343155f
C385 m1_n3334_8532# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.726259f
C386 m1_n3208_8640# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.418123f
C387 m1_18790_1436# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 4.56003f
C388 m1_282_n2232# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.426502f
C389 m1_n3561_8311# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 4.231357f
C390 ibias sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 3.444569f
C391 m1_n3955_n943# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 17.720417f
C392 vb3 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 38.239674f
C393 m1_n5906_n318# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 11.850327f
C394 m1_23556_n2064# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 4.200093f
C395 m1_22524_n1868# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 5.222614f
C396 m1_n5912_464# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 45.838978f
C397 m1_n3667_4379# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.958798f
C398 m1_16202_3432# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 84.157875f
C399 m1_32854_1648# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.101934p
C400 m1_32714_1904# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 98.04854f
C401 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_18/a_50_n200# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.164663f
C402 m1_25484_9858# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.400907f
C403 m1_23420_9858# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.898371f
C404 m1_2256_n728# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 4.89539f
C405 m1_32616_n282# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.558119f
C406 m1_32494_n358# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.724822f
C407 m1_32372_1542# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.557135f
C408 m1_32250_1542# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.720425f
C409 m1_32128_n282# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.55425f
C410 m1_32006_n358# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.706989f
C411 m1_n5902_n1890# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 14.907709f
C412 m1_n4694_n312# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 53.079594f
C413 m1_12142_11768# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.349232f
C414 sky130_fd_pr__nfet_g5v0d10v5_CTEUHA_14/a_50_n200# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.181944f
C415 m1_n3080_8896# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 7.500638f
C416 m1_n3947_7845# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 12.208119f
C417 m1_180_4838# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 8.941923f
C418 m1_790_6356# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 15.466468f
C419 m1_n5902_n1100# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 29.14309f
C420 m1_806_3964# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 10.143394f
C421 m1_180_3630# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 13.001485f
C422 vinp sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 23.89074f
C423 m1_n5904_n2678# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 15.705387f
C424 m1_n5910_1250# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 31.921715f
C425 li_9924_630# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 17.232986f
C426 vinn sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 18.434546f
C427 m1_3549_9621# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.004346f
C428 vout sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 22.613409f
C429 m1_13086_11886# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.614825f
C430 net12 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 8.696936f
C431 m1_n6000_2704# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 12.965477f
C432 m1_779_5148# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 8.414129f
C433 m1_18668_3467# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.185009f
C434 ena sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.227673f
C435 dvdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 3.974578f
C436 m1_791_7588# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 4.63843f
C437 m1_n4698_n3450# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 19.63964f
C438 avdd sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 5.981224p
C439 m1_n2158_9110# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 15.992849f
C440 m1_n4182_7627# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 0.69899f
C441 m1_n3777_8065# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 6.399398f
C442 m1_n4704_472# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 14.688632f
C443 m1_n592_3104# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 25.813177f
C444 m1_n1154_3624# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 12.968743f
C445 net28 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 2.85025f
C446 net29 sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.2079f
C447 m1_n4692_n1074# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 43.43436f
C448 m1_n3264_4838# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 2.542089f
C449 m1_n9267_3854# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 5.232735f
C450 m1_n8442_3847# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 3.812793f
C451 m1_n1846_3922# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 1.660667f
C452 m1_n4685_n1863# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 3.865835f
C453 m1_n3750_n668# sky130_fd_pr__pfet_g5v0d10v5_CVG6CD_13/0 2.094447f
.ends


magic
tech sky130A
magscale 1 2
timestamp 1713232886
<< pwell >>
rect -3553 -708 3553 708
<< mvnmos >>
rect -3325 -450 -3125 450
rect -3067 -450 -2867 450
rect -2809 -450 -2609 450
rect -2551 -450 -2351 450
rect -2293 -450 -2093 450
rect -2035 -450 -1835 450
rect -1777 -450 -1577 450
rect -1519 -450 -1319 450
rect -1261 -450 -1061 450
rect -1003 -450 -803 450
rect -745 -450 -545 450
rect -487 -450 -287 450
rect -229 -450 -29 450
rect 29 -450 229 450
rect 287 -450 487 450
rect 545 -450 745 450
rect 803 -450 1003 450
rect 1061 -450 1261 450
rect 1319 -450 1519 450
rect 1577 -450 1777 450
rect 1835 -450 2035 450
rect 2093 -450 2293 450
rect 2351 -450 2551 450
rect 2609 -450 2809 450
rect 2867 -450 3067 450
rect 3125 -450 3325 450
<< mvndiff >>
rect -3383 438 -3325 450
rect -3383 -438 -3371 438
rect -3337 -438 -3325 438
rect -3383 -450 -3325 -438
rect -3125 438 -3067 450
rect -3125 -438 -3113 438
rect -3079 -438 -3067 438
rect -3125 -450 -3067 -438
rect -2867 438 -2809 450
rect -2867 -438 -2855 438
rect -2821 -438 -2809 438
rect -2867 -450 -2809 -438
rect -2609 438 -2551 450
rect -2609 -438 -2597 438
rect -2563 -438 -2551 438
rect -2609 -450 -2551 -438
rect -2351 438 -2293 450
rect -2351 -438 -2339 438
rect -2305 -438 -2293 438
rect -2351 -450 -2293 -438
rect -2093 438 -2035 450
rect -2093 -438 -2081 438
rect -2047 -438 -2035 438
rect -2093 -450 -2035 -438
rect -1835 438 -1777 450
rect -1835 -438 -1823 438
rect -1789 -438 -1777 438
rect -1835 -450 -1777 -438
rect -1577 438 -1519 450
rect -1577 -438 -1565 438
rect -1531 -438 -1519 438
rect -1577 -450 -1519 -438
rect -1319 438 -1261 450
rect -1319 -438 -1307 438
rect -1273 -438 -1261 438
rect -1319 -450 -1261 -438
rect -1061 438 -1003 450
rect -1061 -438 -1049 438
rect -1015 -438 -1003 438
rect -1061 -450 -1003 -438
rect -803 438 -745 450
rect -803 -438 -791 438
rect -757 -438 -745 438
rect -803 -450 -745 -438
rect -545 438 -487 450
rect -545 -438 -533 438
rect -499 -438 -487 438
rect -545 -450 -487 -438
rect -287 438 -229 450
rect -287 -438 -275 438
rect -241 -438 -229 438
rect -287 -450 -229 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 229 438 287 450
rect 229 -438 241 438
rect 275 -438 287 438
rect 229 -450 287 -438
rect 487 438 545 450
rect 487 -438 499 438
rect 533 -438 545 438
rect 487 -450 545 -438
rect 745 438 803 450
rect 745 -438 757 438
rect 791 -438 803 438
rect 745 -450 803 -438
rect 1003 438 1061 450
rect 1003 -438 1015 438
rect 1049 -438 1061 438
rect 1003 -450 1061 -438
rect 1261 438 1319 450
rect 1261 -438 1273 438
rect 1307 -438 1319 438
rect 1261 -450 1319 -438
rect 1519 438 1577 450
rect 1519 -438 1531 438
rect 1565 -438 1577 438
rect 1519 -450 1577 -438
rect 1777 438 1835 450
rect 1777 -438 1789 438
rect 1823 -438 1835 438
rect 1777 -450 1835 -438
rect 2035 438 2093 450
rect 2035 -438 2047 438
rect 2081 -438 2093 438
rect 2035 -450 2093 -438
rect 2293 438 2351 450
rect 2293 -438 2305 438
rect 2339 -438 2351 438
rect 2293 -450 2351 -438
rect 2551 438 2609 450
rect 2551 -438 2563 438
rect 2597 -438 2609 438
rect 2551 -450 2609 -438
rect 2809 438 2867 450
rect 2809 -438 2821 438
rect 2855 -438 2867 438
rect 2809 -450 2867 -438
rect 3067 438 3125 450
rect 3067 -438 3079 438
rect 3113 -438 3125 438
rect 3067 -450 3125 -438
rect 3325 438 3383 450
rect 3325 -438 3337 438
rect 3371 -438 3383 438
rect 3325 -450 3383 -438
<< mvndiffc >>
rect -3371 -438 -3337 438
rect -3113 -438 -3079 438
rect -2855 -438 -2821 438
rect -2597 -438 -2563 438
rect -2339 -438 -2305 438
rect -2081 -438 -2047 438
rect -1823 -438 -1789 438
rect -1565 -438 -1531 438
rect -1307 -438 -1273 438
rect -1049 -438 -1015 438
rect -791 -438 -757 438
rect -533 -438 -499 438
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
rect 499 -438 533 438
rect 757 -438 791 438
rect 1015 -438 1049 438
rect 1273 -438 1307 438
rect 1531 -438 1565 438
rect 1789 -438 1823 438
rect 2047 -438 2081 438
rect 2305 -438 2339 438
rect 2563 -438 2597 438
rect 2821 -438 2855 438
rect 3079 -438 3113 438
rect 3337 -438 3371 438
<< mvpsubdiff >>
rect -3517 660 3517 672
rect -3517 626 -3409 660
rect 3409 626 3517 660
rect -3517 614 3517 626
rect -3517 564 -3459 614
rect -3517 -564 -3505 564
rect -3471 -564 -3459 564
rect 3459 564 3517 614
rect -3517 -614 -3459 -564
rect 3459 -564 3471 564
rect 3505 -564 3517 564
rect 3459 -614 3517 -564
rect -3517 -626 3517 -614
rect -3517 -660 -3409 -626
rect 3409 -660 3517 -626
rect -3517 -672 3517 -660
<< mvpsubdiffcont >>
rect -3409 626 3409 660
rect -3505 -564 -3471 564
rect 3471 -564 3505 564
rect -3409 -660 3409 -626
<< poly >>
rect -3325 522 -3125 538
rect -3325 488 -3309 522
rect -3141 488 -3125 522
rect -3325 450 -3125 488
rect -3067 522 -2867 538
rect -3067 488 -3051 522
rect -2883 488 -2867 522
rect -3067 450 -2867 488
rect -2809 522 -2609 538
rect -2809 488 -2793 522
rect -2625 488 -2609 522
rect -2809 450 -2609 488
rect -2551 522 -2351 538
rect -2551 488 -2535 522
rect -2367 488 -2351 522
rect -2551 450 -2351 488
rect -2293 522 -2093 538
rect -2293 488 -2277 522
rect -2109 488 -2093 522
rect -2293 450 -2093 488
rect -2035 522 -1835 538
rect -2035 488 -2019 522
rect -1851 488 -1835 522
rect -2035 450 -1835 488
rect -1777 522 -1577 538
rect -1777 488 -1761 522
rect -1593 488 -1577 522
rect -1777 450 -1577 488
rect -1519 522 -1319 538
rect -1519 488 -1503 522
rect -1335 488 -1319 522
rect -1519 450 -1319 488
rect -1261 522 -1061 538
rect -1261 488 -1245 522
rect -1077 488 -1061 522
rect -1261 450 -1061 488
rect -1003 522 -803 538
rect -1003 488 -987 522
rect -819 488 -803 522
rect -1003 450 -803 488
rect -745 522 -545 538
rect -745 488 -729 522
rect -561 488 -545 522
rect -745 450 -545 488
rect -487 522 -287 538
rect -487 488 -471 522
rect -303 488 -287 522
rect -487 450 -287 488
rect -229 522 -29 538
rect -229 488 -213 522
rect -45 488 -29 522
rect -229 450 -29 488
rect 29 522 229 538
rect 29 488 45 522
rect 213 488 229 522
rect 29 450 229 488
rect 287 522 487 538
rect 287 488 303 522
rect 471 488 487 522
rect 287 450 487 488
rect 545 522 745 538
rect 545 488 561 522
rect 729 488 745 522
rect 545 450 745 488
rect 803 522 1003 538
rect 803 488 819 522
rect 987 488 1003 522
rect 803 450 1003 488
rect 1061 522 1261 538
rect 1061 488 1077 522
rect 1245 488 1261 522
rect 1061 450 1261 488
rect 1319 522 1519 538
rect 1319 488 1335 522
rect 1503 488 1519 522
rect 1319 450 1519 488
rect 1577 522 1777 538
rect 1577 488 1593 522
rect 1761 488 1777 522
rect 1577 450 1777 488
rect 1835 522 2035 538
rect 1835 488 1851 522
rect 2019 488 2035 522
rect 1835 450 2035 488
rect 2093 522 2293 538
rect 2093 488 2109 522
rect 2277 488 2293 522
rect 2093 450 2293 488
rect 2351 522 2551 538
rect 2351 488 2367 522
rect 2535 488 2551 522
rect 2351 450 2551 488
rect 2609 522 2809 538
rect 2609 488 2625 522
rect 2793 488 2809 522
rect 2609 450 2809 488
rect 2867 522 3067 538
rect 2867 488 2883 522
rect 3051 488 3067 522
rect 2867 450 3067 488
rect 3125 522 3325 538
rect 3125 488 3141 522
rect 3309 488 3325 522
rect 3125 450 3325 488
rect -3325 -488 -3125 -450
rect -3325 -522 -3309 -488
rect -3141 -522 -3125 -488
rect -3325 -538 -3125 -522
rect -3067 -488 -2867 -450
rect -3067 -522 -3051 -488
rect -2883 -522 -2867 -488
rect -3067 -538 -2867 -522
rect -2809 -488 -2609 -450
rect -2809 -522 -2793 -488
rect -2625 -522 -2609 -488
rect -2809 -538 -2609 -522
rect -2551 -488 -2351 -450
rect -2551 -522 -2535 -488
rect -2367 -522 -2351 -488
rect -2551 -538 -2351 -522
rect -2293 -488 -2093 -450
rect -2293 -522 -2277 -488
rect -2109 -522 -2093 -488
rect -2293 -538 -2093 -522
rect -2035 -488 -1835 -450
rect -2035 -522 -2019 -488
rect -1851 -522 -1835 -488
rect -2035 -538 -1835 -522
rect -1777 -488 -1577 -450
rect -1777 -522 -1761 -488
rect -1593 -522 -1577 -488
rect -1777 -538 -1577 -522
rect -1519 -488 -1319 -450
rect -1519 -522 -1503 -488
rect -1335 -522 -1319 -488
rect -1519 -538 -1319 -522
rect -1261 -488 -1061 -450
rect -1261 -522 -1245 -488
rect -1077 -522 -1061 -488
rect -1261 -538 -1061 -522
rect -1003 -488 -803 -450
rect -1003 -522 -987 -488
rect -819 -522 -803 -488
rect -1003 -538 -803 -522
rect -745 -488 -545 -450
rect -745 -522 -729 -488
rect -561 -522 -545 -488
rect -745 -538 -545 -522
rect -487 -488 -287 -450
rect -487 -522 -471 -488
rect -303 -522 -287 -488
rect -487 -538 -287 -522
rect -229 -488 -29 -450
rect -229 -522 -213 -488
rect -45 -522 -29 -488
rect -229 -538 -29 -522
rect 29 -488 229 -450
rect 29 -522 45 -488
rect 213 -522 229 -488
rect 29 -538 229 -522
rect 287 -488 487 -450
rect 287 -522 303 -488
rect 471 -522 487 -488
rect 287 -538 487 -522
rect 545 -488 745 -450
rect 545 -522 561 -488
rect 729 -522 745 -488
rect 545 -538 745 -522
rect 803 -488 1003 -450
rect 803 -522 819 -488
rect 987 -522 1003 -488
rect 803 -538 1003 -522
rect 1061 -488 1261 -450
rect 1061 -522 1077 -488
rect 1245 -522 1261 -488
rect 1061 -538 1261 -522
rect 1319 -488 1519 -450
rect 1319 -522 1335 -488
rect 1503 -522 1519 -488
rect 1319 -538 1519 -522
rect 1577 -488 1777 -450
rect 1577 -522 1593 -488
rect 1761 -522 1777 -488
rect 1577 -538 1777 -522
rect 1835 -488 2035 -450
rect 1835 -522 1851 -488
rect 2019 -522 2035 -488
rect 1835 -538 2035 -522
rect 2093 -488 2293 -450
rect 2093 -522 2109 -488
rect 2277 -522 2293 -488
rect 2093 -538 2293 -522
rect 2351 -488 2551 -450
rect 2351 -522 2367 -488
rect 2535 -522 2551 -488
rect 2351 -538 2551 -522
rect 2609 -488 2809 -450
rect 2609 -522 2625 -488
rect 2793 -522 2809 -488
rect 2609 -538 2809 -522
rect 2867 -488 3067 -450
rect 2867 -522 2883 -488
rect 3051 -522 3067 -488
rect 2867 -538 3067 -522
rect 3125 -488 3325 -450
rect 3125 -522 3141 -488
rect 3309 -522 3325 -488
rect 3125 -538 3325 -522
<< polycont >>
rect -3309 488 -3141 522
rect -3051 488 -2883 522
rect -2793 488 -2625 522
rect -2535 488 -2367 522
rect -2277 488 -2109 522
rect -2019 488 -1851 522
rect -1761 488 -1593 522
rect -1503 488 -1335 522
rect -1245 488 -1077 522
rect -987 488 -819 522
rect -729 488 -561 522
rect -471 488 -303 522
rect -213 488 -45 522
rect 45 488 213 522
rect 303 488 471 522
rect 561 488 729 522
rect 819 488 987 522
rect 1077 488 1245 522
rect 1335 488 1503 522
rect 1593 488 1761 522
rect 1851 488 2019 522
rect 2109 488 2277 522
rect 2367 488 2535 522
rect 2625 488 2793 522
rect 2883 488 3051 522
rect 3141 488 3309 522
rect -3309 -522 -3141 -488
rect -3051 -522 -2883 -488
rect -2793 -522 -2625 -488
rect -2535 -522 -2367 -488
rect -2277 -522 -2109 -488
rect -2019 -522 -1851 -488
rect -1761 -522 -1593 -488
rect -1503 -522 -1335 -488
rect -1245 -522 -1077 -488
rect -987 -522 -819 -488
rect -729 -522 -561 -488
rect -471 -522 -303 -488
rect -213 -522 -45 -488
rect 45 -522 213 -488
rect 303 -522 471 -488
rect 561 -522 729 -488
rect 819 -522 987 -488
rect 1077 -522 1245 -488
rect 1335 -522 1503 -488
rect 1593 -522 1761 -488
rect 1851 -522 2019 -488
rect 2109 -522 2277 -488
rect 2367 -522 2535 -488
rect 2625 -522 2793 -488
rect 2883 -522 3051 -488
rect 3141 -522 3309 -488
<< locali >>
rect -3505 626 -3409 660
rect 3409 626 3505 660
rect -3505 564 -3471 626
rect 3471 564 3505 626
rect -3325 488 -3309 522
rect -3141 488 -3125 522
rect -3067 488 -3051 522
rect -2883 488 -2867 522
rect -2809 488 -2793 522
rect -2625 488 -2609 522
rect -2551 488 -2535 522
rect -2367 488 -2351 522
rect -2293 488 -2277 522
rect -2109 488 -2093 522
rect -2035 488 -2019 522
rect -1851 488 -1835 522
rect -1777 488 -1761 522
rect -1593 488 -1577 522
rect -1519 488 -1503 522
rect -1335 488 -1319 522
rect -1261 488 -1245 522
rect -1077 488 -1061 522
rect -1003 488 -987 522
rect -819 488 -803 522
rect -745 488 -729 522
rect -561 488 -545 522
rect -487 488 -471 522
rect -303 488 -287 522
rect -229 488 -213 522
rect -45 488 -29 522
rect 29 488 45 522
rect 213 488 229 522
rect 287 488 303 522
rect 471 488 487 522
rect 545 488 561 522
rect 729 488 745 522
rect 803 488 819 522
rect 987 488 1003 522
rect 1061 488 1077 522
rect 1245 488 1261 522
rect 1319 488 1335 522
rect 1503 488 1519 522
rect 1577 488 1593 522
rect 1761 488 1777 522
rect 1835 488 1851 522
rect 2019 488 2035 522
rect 2093 488 2109 522
rect 2277 488 2293 522
rect 2351 488 2367 522
rect 2535 488 2551 522
rect 2609 488 2625 522
rect 2793 488 2809 522
rect 2867 488 2883 522
rect 3051 488 3067 522
rect 3125 488 3141 522
rect 3309 488 3325 522
rect -3371 438 -3337 454
rect -3371 -454 -3337 -438
rect -3113 438 -3079 454
rect -3113 -454 -3079 -438
rect -2855 438 -2821 454
rect -2855 -454 -2821 -438
rect -2597 438 -2563 454
rect -2597 -454 -2563 -438
rect -2339 438 -2305 454
rect -2339 -454 -2305 -438
rect -2081 438 -2047 454
rect -2081 -454 -2047 -438
rect -1823 438 -1789 454
rect -1823 -454 -1789 -438
rect -1565 438 -1531 454
rect -1565 -454 -1531 -438
rect -1307 438 -1273 454
rect -1307 -454 -1273 -438
rect -1049 438 -1015 454
rect -1049 -454 -1015 -438
rect -791 438 -757 454
rect -791 -454 -757 -438
rect -533 438 -499 454
rect -533 -454 -499 -438
rect -275 438 -241 454
rect -275 -454 -241 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 241 438 275 454
rect 241 -454 275 -438
rect 499 438 533 454
rect 499 -454 533 -438
rect 757 438 791 454
rect 757 -454 791 -438
rect 1015 438 1049 454
rect 1015 -454 1049 -438
rect 1273 438 1307 454
rect 1273 -454 1307 -438
rect 1531 438 1565 454
rect 1531 -454 1565 -438
rect 1789 438 1823 454
rect 1789 -454 1823 -438
rect 2047 438 2081 454
rect 2047 -454 2081 -438
rect 2305 438 2339 454
rect 2305 -454 2339 -438
rect 2563 438 2597 454
rect 2563 -454 2597 -438
rect 2821 438 2855 454
rect 2821 -454 2855 -438
rect 3079 438 3113 454
rect 3079 -454 3113 -438
rect 3337 438 3371 454
rect 3337 -454 3371 -438
rect -3325 -522 -3309 -488
rect -3141 -522 -3125 -488
rect -3067 -522 -3051 -488
rect -2883 -522 -2867 -488
rect -2809 -522 -2793 -488
rect -2625 -522 -2609 -488
rect -2551 -522 -2535 -488
rect -2367 -522 -2351 -488
rect -2293 -522 -2277 -488
rect -2109 -522 -2093 -488
rect -2035 -522 -2019 -488
rect -1851 -522 -1835 -488
rect -1777 -522 -1761 -488
rect -1593 -522 -1577 -488
rect -1519 -522 -1503 -488
rect -1335 -522 -1319 -488
rect -1261 -522 -1245 -488
rect -1077 -522 -1061 -488
rect -1003 -522 -987 -488
rect -819 -522 -803 -488
rect -745 -522 -729 -488
rect -561 -522 -545 -488
rect -487 -522 -471 -488
rect -303 -522 -287 -488
rect -229 -522 -213 -488
rect -45 -522 -29 -488
rect 29 -522 45 -488
rect 213 -522 229 -488
rect 287 -522 303 -488
rect 471 -522 487 -488
rect 545 -522 561 -488
rect 729 -522 745 -488
rect 803 -522 819 -488
rect 987 -522 1003 -488
rect 1061 -522 1077 -488
rect 1245 -522 1261 -488
rect 1319 -522 1335 -488
rect 1503 -522 1519 -488
rect 1577 -522 1593 -488
rect 1761 -522 1777 -488
rect 1835 -522 1851 -488
rect 2019 -522 2035 -488
rect 2093 -522 2109 -488
rect 2277 -522 2293 -488
rect 2351 -522 2367 -488
rect 2535 -522 2551 -488
rect 2609 -522 2625 -488
rect 2793 -522 2809 -488
rect 2867 -522 2883 -488
rect 3051 -522 3067 -488
rect 3125 -522 3141 -488
rect 3309 -522 3325 -488
rect -3505 -626 -3471 -564
rect 3471 -626 3505 -564
rect -3505 -660 -3409 -626
rect 3409 -660 3505 -626
<< viali >>
rect -3309 488 -3141 522
rect -3051 488 -2883 522
rect -2793 488 -2625 522
rect -2535 488 -2367 522
rect -2277 488 -2109 522
rect -2019 488 -1851 522
rect -1761 488 -1593 522
rect -1503 488 -1335 522
rect -1245 488 -1077 522
rect -987 488 -819 522
rect -729 488 -561 522
rect -471 488 -303 522
rect -213 488 -45 522
rect 45 488 213 522
rect 303 488 471 522
rect 561 488 729 522
rect 819 488 987 522
rect 1077 488 1245 522
rect 1335 488 1503 522
rect 1593 488 1761 522
rect 1851 488 2019 522
rect 2109 488 2277 522
rect 2367 488 2535 522
rect 2625 488 2793 522
rect 2883 488 3051 522
rect 3141 488 3309 522
rect -3371 -438 -3337 438
rect -3113 -438 -3079 438
rect -2855 -438 -2821 438
rect -2597 -438 -2563 438
rect -2339 -438 -2305 438
rect -2081 -438 -2047 438
rect -1823 -438 -1789 438
rect -1565 -438 -1531 438
rect -1307 -438 -1273 438
rect -1049 -438 -1015 438
rect -791 -438 -757 438
rect -533 -438 -499 438
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
rect 499 -438 533 438
rect 757 -438 791 438
rect 1015 -438 1049 438
rect 1273 -438 1307 438
rect 1531 -438 1565 438
rect 1789 -438 1823 438
rect 2047 -438 2081 438
rect 2305 -438 2339 438
rect 2563 -438 2597 438
rect 2821 -438 2855 438
rect 3079 -438 3113 438
rect 3337 -438 3371 438
rect -3309 -522 -3141 -488
rect -3051 -522 -2883 -488
rect -2793 -522 -2625 -488
rect -2535 -522 -2367 -488
rect -2277 -522 -2109 -488
rect -2019 -522 -1851 -488
rect -1761 -522 -1593 -488
rect -1503 -522 -1335 -488
rect -1245 -522 -1077 -488
rect -987 -522 -819 -488
rect -729 -522 -561 -488
rect -471 -522 -303 -488
rect -213 -522 -45 -488
rect 45 -522 213 -488
rect 303 -522 471 -488
rect 561 -522 729 -488
rect 819 -522 987 -488
rect 1077 -522 1245 -488
rect 1335 -522 1503 -488
rect 1593 -522 1761 -488
rect 1851 -522 2019 -488
rect 2109 -522 2277 -488
rect 2367 -522 2535 -488
rect 2625 -522 2793 -488
rect 2883 -522 3051 -488
rect 3141 -522 3309 -488
<< metal1 >>
rect -3321 522 -3129 528
rect -3321 488 -3309 522
rect -3141 488 -3129 522
rect -3321 482 -3129 488
rect -3063 522 -2871 528
rect -3063 488 -3051 522
rect -2883 488 -2871 522
rect -3063 482 -2871 488
rect -2805 522 -2613 528
rect -2805 488 -2793 522
rect -2625 488 -2613 522
rect -2805 482 -2613 488
rect -2547 522 -2355 528
rect -2547 488 -2535 522
rect -2367 488 -2355 522
rect -2547 482 -2355 488
rect -2289 522 -2097 528
rect -2289 488 -2277 522
rect -2109 488 -2097 522
rect -2289 482 -2097 488
rect -2031 522 -1839 528
rect -2031 488 -2019 522
rect -1851 488 -1839 522
rect -2031 482 -1839 488
rect -1773 522 -1581 528
rect -1773 488 -1761 522
rect -1593 488 -1581 522
rect -1773 482 -1581 488
rect -1515 522 -1323 528
rect -1515 488 -1503 522
rect -1335 488 -1323 522
rect -1515 482 -1323 488
rect -1257 522 -1065 528
rect -1257 488 -1245 522
rect -1077 488 -1065 522
rect -1257 482 -1065 488
rect -999 522 -807 528
rect -999 488 -987 522
rect -819 488 -807 522
rect -999 482 -807 488
rect -741 522 -549 528
rect -741 488 -729 522
rect -561 488 -549 522
rect -741 482 -549 488
rect -483 522 -291 528
rect -483 488 -471 522
rect -303 488 -291 522
rect -483 482 -291 488
rect -225 522 -33 528
rect -225 488 -213 522
rect -45 488 -33 522
rect -225 482 -33 488
rect 33 522 225 528
rect 33 488 45 522
rect 213 488 225 522
rect 33 482 225 488
rect 291 522 483 528
rect 291 488 303 522
rect 471 488 483 522
rect 291 482 483 488
rect 549 522 741 528
rect 549 488 561 522
rect 729 488 741 522
rect 549 482 741 488
rect 807 522 999 528
rect 807 488 819 522
rect 987 488 999 522
rect 807 482 999 488
rect 1065 522 1257 528
rect 1065 488 1077 522
rect 1245 488 1257 522
rect 1065 482 1257 488
rect 1323 522 1515 528
rect 1323 488 1335 522
rect 1503 488 1515 522
rect 1323 482 1515 488
rect 1581 522 1773 528
rect 1581 488 1593 522
rect 1761 488 1773 522
rect 1581 482 1773 488
rect 1839 522 2031 528
rect 1839 488 1851 522
rect 2019 488 2031 522
rect 1839 482 2031 488
rect 2097 522 2289 528
rect 2097 488 2109 522
rect 2277 488 2289 522
rect 2097 482 2289 488
rect 2355 522 2547 528
rect 2355 488 2367 522
rect 2535 488 2547 522
rect 2355 482 2547 488
rect 2613 522 2805 528
rect 2613 488 2625 522
rect 2793 488 2805 522
rect 2613 482 2805 488
rect 2871 522 3063 528
rect 2871 488 2883 522
rect 3051 488 3063 522
rect 2871 482 3063 488
rect 3129 522 3321 528
rect 3129 488 3141 522
rect 3309 488 3321 522
rect 3129 482 3321 488
rect -3377 438 -3331 450
rect -3377 -438 -3371 438
rect -3337 -438 -3331 438
rect -3377 -450 -3331 -438
rect -3119 438 -3073 450
rect -3119 -438 -3113 438
rect -3079 -438 -3073 438
rect -3119 -450 -3073 -438
rect -2861 438 -2815 450
rect -2861 -438 -2855 438
rect -2821 -438 -2815 438
rect -2861 -450 -2815 -438
rect -2603 438 -2557 450
rect -2603 -438 -2597 438
rect -2563 -438 -2557 438
rect -2603 -450 -2557 -438
rect -2345 438 -2299 450
rect -2345 -438 -2339 438
rect -2305 -438 -2299 438
rect -2345 -450 -2299 -438
rect -2087 438 -2041 450
rect -2087 -438 -2081 438
rect -2047 -438 -2041 438
rect -2087 -450 -2041 -438
rect -1829 438 -1783 450
rect -1829 -438 -1823 438
rect -1789 -438 -1783 438
rect -1829 -450 -1783 -438
rect -1571 438 -1525 450
rect -1571 -438 -1565 438
rect -1531 -438 -1525 438
rect -1571 -450 -1525 -438
rect -1313 438 -1267 450
rect -1313 -438 -1307 438
rect -1273 -438 -1267 438
rect -1313 -450 -1267 -438
rect -1055 438 -1009 450
rect -1055 -438 -1049 438
rect -1015 -438 -1009 438
rect -1055 -450 -1009 -438
rect -797 438 -751 450
rect -797 -438 -791 438
rect -757 -438 -751 438
rect -797 -450 -751 -438
rect -539 438 -493 450
rect -539 -438 -533 438
rect -499 -438 -493 438
rect -539 -450 -493 -438
rect -281 438 -235 450
rect -281 -438 -275 438
rect -241 -438 -235 438
rect -281 -450 -235 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 235 438 281 450
rect 235 -438 241 438
rect 275 -438 281 438
rect 235 -450 281 -438
rect 493 438 539 450
rect 493 -438 499 438
rect 533 -438 539 438
rect 493 -450 539 -438
rect 751 438 797 450
rect 751 -438 757 438
rect 791 -438 797 438
rect 751 -450 797 -438
rect 1009 438 1055 450
rect 1009 -438 1015 438
rect 1049 -438 1055 438
rect 1009 -450 1055 -438
rect 1267 438 1313 450
rect 1267 -438 1273 438
rect 1307 -438 1313 438
rect 1267 -450 1313 -438
rect 1525 438 1571 450
rect 1525 -438 1531 438
rect 1565 -438 1571 438
rect 1525 -450 1571 -438
rect 1783 438 1829 450
rect 1783 -438 1789 438
rect 1823 -438 1829 438
rect 1783 -450 1829 -438
rect 2041 438 2087 450
rect 2041 -438 2047 438
rect 2081 -438 2087 438
rect 2041 -450 2087 -438
rect 2299 438 2345 450
rect 2299 -438 2305 438
rect 2339 -438 2345 438
rect 2299 -450 2345 -438
rect 2557 438 2603 450
rect 2557 -438 2563 438
rect 2597 -438 2603 438
rect 2557 -450 2603 -438
rect 2815 438 2861 450
rect 2815 -438 2821 438
rect 2855 -438 2861 438
rect 2815 -450 2861 -438
rect 3073 438 3119 450
rect 3073 -438 3079 438
rect 3113 -438 3119 438
rect 3073 -450 3119 -438
rect 3331 438 3377 450
rect 3331 -438 3337 438
rect 3371 -438 3377 438
rect 3331 -450 3377 -438
rect -3321 -488 -3129 -482
rect -3321 -522 -3309 -488
rect -3141 -522 -3129 -488
rect -3321 -528 -3129 -522
rect -3063 -488 -2871 -482
rect -3063 -522 -3051 -488
rect -2883 -522 -2871 -488
rect -3063 -528 -2871 -522
rect -2805 -488 -2613 -482
rect -2805 -522 -2793 -488
rect -2625 -522 -2613 -488
rect -2805 -528 -2613 -522
rect -2547 -488 -2355 -482
rect -2547 -522 -2535 -488
rect -2367 -522 -2355 -488
rect -2547 -528 -2355 -522
rect -2289 -488 -2097 -482
rect -2289 -522 -2277 -488
rect -2109 -522 -2097 -488
rect -2289 -528 -2097 -522
rect -2031 -488 -1839 -482
rect -2031 -522 -2019 -488
rect -1851 -522 -1839 -488
rect -2031 -528 -1839 -522
rect -1773 -488 -1581 -482
rect -1773 -522 -1761 -488
rect -1593 -522 -1581 -488
rect -1773 -528 -1581 -522
rect -1515 -488 -1323 -482
rect -1515 -522 -1503 -488
rect -1335 -522 -1323 -488
rect -1515 -528 -1323 -522
rect -1257 -488 -1065 -482
rect -1257 -522 -1245 -488
rect -1077 -522 -1065 -488
rect -1257 -528 -1065 -522
rect -999 -488 -807 -482
rect -999 -522 -987 -488
rect -819 -522 -807 -488
rect -999 -528 -807 -522
rect -741 -488 -549 -482
rect -741 -522 -729 -488
rect -561 -522 -549 -488
rect -741 -528 -549 -522
rect -483 -488 -291 -482
rect -483 -522 -471 -488
rect -303 -522 -291 -488
rect -483 -528 -291 -522
rect -225 -488 -33 -482
rect -225 -522 -213 -488
rect -45 -522 -33 -488
rect -225 -528 -33 -522
rect 33 -488 225 -482
rect 33 -522 45 -488
rect 213 -522 225 -488
rect 33 -528 225 -522
rect 291 -488 483 -482
rect 291 -522 303 -488
rect 471 -522 483 -488
rect 291 -528 483 -522
rect 549 -488 741 -482
rect 549 -522 561 -488
rect 729 -522 741 -488
rect 549 -528 741 -522
rect 807 -488 999 -482
rect 807 -522 819 -488
rect 987 -522 999 -488
rect 807 -528 999 -522
rect 1065 -488 1257 -482
rect 1065 -522 1077 -488
rect 1245 -522 1257 -488
rect 1065 -528 1257 -522
rect 1323 -488 1515 -482
rect 1323 -522 1335 -488
rect 1503 -522 1515 -488
rect 1323 -528 1515 -522
rect 1581 -488 1773 -482
rect 1581 -522 1593 -488
rect 1761 -522 1773 -488
rect 1581 -528 1773 -522
rect 1839 -488 2031 -482
rect 1839 -522 1851 -488
rect 2019 -522 2031 -488
rect 1839 -528 2031 -522
rect 2097 -488 2289 -482
rect 2097 -522 2109 -488
rect 2277 -522 2289 -488
rect 2097 -528 2289 -522
rect 2355 -488 2547 -482
rect 2355 -522 2367 -488
rect 2535 -522 2547 -488
rect 2355 -528 2547 -522
rect 2613 -488 2805 -482
rect 2613 -522 2625 -488
rect 2793 -522 2805 -488
rect 2613 -528 2805 -522
rect 2871 -488 3063 -482
rect 2871 -522 2883 -488
rect 3051 -522 3063 -488
rect 2871 -528 3063 -522
rect 3129 -488 3321 -482
rect 3129 -522 3141 -488
rect 3309 -522 3321 -488
rect 3129 -528 3321 -522
<< properties >>
string FIXED_BBOX -3488 -643 3488 643
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 1 m 1 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

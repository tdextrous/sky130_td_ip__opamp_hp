magic
tech sky130A
magscale 1 2
timestamp 1713391144
<< nwell >>
rect -4615 -2797 4615 2797
<< mvpmos >>
rect -4357 -2500 -4157 2500
rect -4099 -2500 -3899 2500
rect -3841 -2500 -3641 2500
rect -3583 -2500 -3383 2500
rect -3325 -2500 -3125 2500
rect -3067 -2500 -2867 2500
rect -2809 -2500 -2609 2500
rect -2551 -2500 -2351 2500
rect -2293 -2500 -2093 2500
rect -2035 -2500 -1835 2500
rect -1777 -2500 -1577 2500
rect -1519 -2500 -1319 2500
rect -1261 -2500 -1061 2500
rect -1003 -2500 -803 2500
rect -745 -2500 -545 2500
rect -487 -2500 -287 2500
rect -229 -2500 -29 2500
rect 29 -2500 229 2500
rect 287 -2500 487 2500
rect 545 -2500 745 2500
rect 803 -2500 1003 2500
rect 1061 -2500 1261 2500
rect 1319 -2500 1519 2500
rect 1577 -2500 1777 2500
rect 1835 -2500 2035 2500
rect 2093 -2500 2293 2500
rect 2351 -2500 2551 2500
rect 2609 -2500 2809 2500
rect 2867 -2500 3067 2500
rect 3125 -2500 3325 2500
rect 3383 -2500 3583 2500
rect 3641 -2500 3841 2500
rect 3899 -2500 4099 2500
rect 4157 -2500 4357 2500
<< mvpdiff >>
rect -4415 2488 -4357 2500
rect -4415 -2488 -4403 2488
rect -4369 -2488 -4357 2488
rect -4415 -2500 -4357 -2488
rect -4157 2488 -4099 2500
rect -4157 -2488 -4145 2488
rect -4111 -2488 -4099 2488
rect -4157 -2500 -4099 -2488
rect -3899 2488 -3841 2500
rect -3899 -2488 -3887 2488
rect -3853 -2488 -3841 2488
rect -3899 -2500 -3841 -2488
rect -3641 2488 -3583 2500
rect -3641 -2488 -3629 2488
rect -3595 -2488 -3583 2488
rect -3641 -2500 -3583 -2488
rect -3383 2488 -3325 2500
rect -3383 -2488 -3371 2488
rect -3337 -2488 -3325 2488
rect -3383 -2500 -3325 -2488
rect -3125 2488 -3067 2500
rect -3125 -2488 -3113 2488
rect -3079 -2488 -3067 2488
rect -3125 -2500 -3067 -2488
rect -2867 2488 -2809 2500
rect -2867 -2488 -2855 2488
rect -2821 -2488 -2809 2488
rect -2867 -2500 -2809 -2488
rect -2609 2488 -2551 2500
rect -2609 -2488 -2597 2488
rect -2563 -2488 -2551 2488
rect -2609 -2500 -2551 -2488
rect -2351 2488 -2293 2500
rect -2351 -2488 -2339 2488
rect -2305 -2488 -2293 2488
rect -2351 -2500 -2293 -2488
rect -2093 2488 -2035 2500
rect -2093 -2488 -2081 2488
rect -2047 -2488 -2035 2488
rect -2093 -2500 -2035 -2488
rect -1835 2488 -1777 2500
rect -1835 -2488 -1823 2488
rect -1789 -2488 -1777 2488
rect -1835 -2500 -1777 -2488
rect -1577 2488 -1519 2500
rect -1577 -2488 -1565 2488
rect -1531 -2488 -1519 2488
rect -1577 -2500 -1519 -2488
rect -1319 2488 -1261 2500
rect -1319 -2488 -1307 2488
rect -1273 -2488 -1261 2488
rect -1319 -2500 -1261 -2488
rect -1061 2488 -1003 2500
rect -1061 -2488 -1049 2488
rect -1015 -2488 -1003 2488
rect -1061 -2500 -1003 -2488
rect -803 2488 -745 2500
rect -803 -2488 -791 2488
rect -757 -2488 -745 2488
rect -803 -2500 -745 -2488
rect -545 2488 -487 2500
rect -545 -2488 -533 2488
rect -499 -2488 -487 2488
rect -545 -2500 -487 -2488
rect -287 2488 -229 2500
rect -287 -2488 -275 2488
rect -241 -2488 -229 2488
rect -287 -2500 -229 -2488
rect -29 2488 29 2500
rect -29 -2488 -17 2488
rect 17 -2488 29 2488
rect -29 -2500 29 -2488
rect 229 2488 287 2500
rect 229 -2488 241 2488
rect 275 -2488 287 2488
rect 229 -2500 287 -2488
rect 487 2488 545 2500
rect 487 -2488 499 2488
rect 533 -2488 545 2488
rect 487 -2500 545 -2488
rect 745 2488 803 2500
rect 745 -2488 757 2488
rect 791 -2488 803 2488
rect 745 -2500 803 -2488
rect 1003 2488 1061 2500
rect 1003 -2488 1015 2488
rect 1049 -2488 1061 2488
rect 1003 -2500 1061 -2488
rect 1261 2488 1319 2500
rect 1261 -2488 1273 2488
rect 1307 -2488 1319 2488
rect 1261 -2500 1319 -2488
rect 1519 2488 1577 2500
rect 1519 -2488 1531 2488
rect 1565 -2488 1577 2488
rect 1519 -2500 1577 -2488
rect 1777 2488 1835 2500
rect 1777 -2488 1789 2488
rect 1823 -2488 1835 2488
rect 1777 -2500 1835 -2488
rect 2035 2488 2093 2500
rect 2035 -2488 2047 2488
rect 2081 -2488 2093 2488
rect 2035 -2500 2093 -2488
rect 2293 2488 2351 2500
rect 2293 -2488 2305 2488
rect 2339 -2488 2351 2488
rect 2293 -2500 2351 -2488
rect 2551 2488 2609 2500
rect 2551 -2488 2563 2488
rect 2597 -2488 2609 2488
rect 2551 -2500 2609 -2488
rect 2809 2488 2867 2500
rect 2809 -2488 2821 2488
rect 2855 -2488 2867 2488
rect 2809 -2500 2867 -2488
rect 3067 2488 3125 2500
rect 3067 -2488 3079 2488
rect 3113 -2488 3125 2488
rect 3067 -2500 3125 -2488
rect 3325 2488 3383 2500
rect 3325 -2488 3337 2488
rect 3371 -2488 3383 2488
rect 3325 -2500 3383 -2488
rect 3583 2488 3641 2500
rect 3583 -2488 3595 2488
rect 3629 -2488 3641 2488
rect 3583 -2500 3641 -2488
rect 3841 2488 3899 2500
rect 3841 -2488 3853 2488
rect 3887 -2488 3899 2488
rect 3841 -2500 3899 -2488
rect 4099 2488 4157 2500
rect 4099 -2488 4111 2488
rect 4145 -2488 4157 2488
rect 4099 -2500 4157 -2488
rect 4357 2488 4415 2500
rect 4357 -2488 4369 2488
rect 4403 -2488 4415 2488
rect 4357 -2500 4415 -2488
<< mvpdiffc >>
rect -4403 -2488 -4369 2488
rect -4145 -2488 -4111 2488
rect -3887 -2488 -3853 2488
rect -3629 -2488 -3595 2488
rect -3371 -2488 -3337 2488
rect -3113 -2488 -3079 2488
rect -2855 -2488 -2821 2488
rect -2597 -2488 -2563 2488
rect -2339 -2488 -2305 2488
rect -2081 -2488 -2047 2488
rect -1823 -2488 -1789 2488
rect -1565 -2488 -1531 2488
rect -1307 -2488 -1273 2488
rect -1049 -2488 -1015 2488
rect -791 -2488 -757 2488
rect -533 -2488 -499 2488
rect -275 -2488 -241 2488
rect -17 -2488 17 2488
rect 241 -2488 275 2488
rect 499 -2488 533 2488
rect 757 -2488 791 2488
rect 1015 -2488 1049 2488
rect 1273 -2488 1307 2488
rect 1531 -2488 1565 2488
rect 1789 -2488 1823 2488
rect 2047 -2488 2081 2488
rect 2305 -2488 2339 2488
rect 2563 -2488 2597 2488
rect 2821 -2488 2855 2488
rect 3079 -2488 3113 2488
rect 3337 -2488 3371 2488
rect 3595 -2488 3629 2488
rect 3853 -2488 3887 2488
rect 4111 -2488 4145 2488
rect 4369 -2488 4403 2488
<< mvnsubdiff >>
rect -4549 2719 4549 2731
rect -4549 2685 -4441 2719
rect 4441 2685 4549 2719
rect -4549 2673 4549 2685
rect -4549 2623 -4491 2673
rect -4549 -2623 -4537 2623
rect -4503 -2623 -4491 2623
rect 4491 2623 4549 2673
rect -4549 -2673 -4491 -2623
rect 4491 -2623 4503 2623
rect 4537 -2623 4549 2623
rect 4491 -2673 4549 -2623
rect -4549 -2685 4549 -2673
rect -4549 -2719 -4441 -2685
rect 4441 -2719 4549 -2685
rect -4549 -2731 4549 -2719
<< mvnsubdiffcont >>
rect -4441 2685 4441 2719
rect -4537 -2623 -4503 2623
rect 4503 -2623 4537 2623
rect -4441 -2719 4441 -2685
<< poly >>
rect -4323 2581 -4191 2597
rect -4323 2564 -4307 2581
rect -4357 2547 -4307 2564
rect -4207 2564 -4191 2581
rect -4065 2581 -3933 2597
rect -4065 2564 -4049 2581
rect -4207 2547 -4157 2564
rect -4357 2500 -4157 2547
rect -4099 2547 -4049 2564
rect -3949 2564 -3933 2581
rect -3807 2581 -3675 2597
rect -3807 2564 -3791 2581
rect -3949 2547 -3899 2564
rect -4099 2500 -3899 2547
rect -3841 2547 -3791 2564
rect -3691 2564 -3675 2581
rect -3549 2581 -3417 2597
rect -3549 2564 -3533 2581
rect -3691 2547 -3641 2564
rect -3841 2500 -3641 2547
rect -3583 2547 -3533 2564
rect -3433 2564 -3417 2581
rect -3291 2581 -3159 2597
rect -3291 2564 -3275 2581
rect -3433 2547 -3383 2564
rect -3583 2500 -3383 2547
rect -3325 2547 -3275 2564
rect -3175 2564 -3159 2581
rect -3033 2581 -2901 2597
rect -3033 2564 -3017 2581
rect -3175 2547 -3125 2564
rect -3325 2500 -3125 2547
rect -3067 2547 -3017 2564
rect -2917 2564 -2901 2581
rect -2775 2581 -2643 2597
rect -2775 2564 -2759 2581
rect -2917 2547 -2867 2564
rect -3067 2500 -2867 2547
rect -2809 2547 -2759 2564
rect -2659 2564 -2643 2581
rect -2517 2581 -2385 2597
rect -2517 2564 -2501 2581
rect -2659 2547 -2609 2564
rect -2809 2500 -2609 2547
rect -2551 2547 -2501 2564
rect -2401 2564 -2385 2581
rect -2259 2581 -2127 2597
rect -2259 2564 -2243 2581
rect -2401 2547 -2351 2564
rect -2551 2500 -2351 2547
rect -2293 2547 -2243 2564
rect -2143 2564 -2127 2581
rect -2001 2581 -1869 2597
rect -2001 2564 -1985 2581
rect -2143 2547 -2093 2564
rect -2293 2500 -2093 2547
rect -2035 2547 -1985 2564
rect -1885 2564 -1869 2581
rect -1743 2581 -1611 2597
rect -1743 2564 -1727 2581
rect -1885 2547 -1835 2564
rect -2035 2500 -1835 2547
rect -1777 2547 -1727 2564
rect -1627 2564 -1611 2581
rect -1485 2581 -1353 2597
rect -1485 2564 -1469 2581
rect -1627 2547 -1577 2564
rect -1777 2500 -1577 2547
rect -1519 2547 -1469 2564
rect -1369 2564 -1353 2581
rect -1227 2581 -1095 2597
rect -1227 2564 -1211 2581
rect -1369 2547 -1319 2564
rect -1519 2500 -1319 2547
rect -1261 2547 -1211 2564
rect -1111 2564 -1095 2581
rect -969 2581 -837 2597
rect -969 2564 -953 2581
rect -1111 2547 -1061 2564
rect -1261 2500 -1061 2547
rect -1003 2547 -953 2564
rect -853 2564 -837 2581
rect -711 2581 -579 2597
rect -711 2564 -695 2581
rect -853 2547 -803 2564
rect -1003 2500 -803 2547
rect -745 2547 -695 2564
rect -595 2564 -579 2581
rect -453 2581 -321 2597
rect -453 2564 -437 2581
rect -595 2547 -545 2564
rect -745 2500 -545 2547
rect -487 2547 -437 2564
rect -337 2564 -321 2581
rect -195 2581 -63 2597
rect -195 2564 -179 2581
rect -337 2547 -287 2564
rect -487 2500 -287 2547
rect -229 2547 -179 2564
rect -79 2564 -63 2581
rect 63 2581 195 2597
rect 63 2564 79 2581
rect -79 2547 -29 2564
rect -229 2500 -29 2547
rect 29 2547 79 2564
rect 179 2564 195 2581
rect 321 2581 453 2597
rect 321 2564 337 2581
rect 179 2547 229 2564
rect 29 2500 229 2547
rect 287 2547 337 2564
rect 437 2564 453 2581
rect 579 2581 711 2597
rect 579 2564 595 2581
rect 437 2547 487 2564
rect 287 2500 487 2547
rect 545 2547 595 2564
rect 695 2564 711 2581
rect 837 2581 969 2597
rect 837 2564 853 2581
rect 695 2547 745 2564
rect 545 2500 745 2547
rect 803 2547 853 2564
rect 953 2564 969 2581
rect 1095 2581 1227 2597
rect 1095 2564 1111 2581
rect 953 2547 1003 2564
rect 803 2500 1003 2547
rect 1061 2547 1111 2564
rect 1211 2564 1227 2581
rect 1353 2581 1485 2597
rect 1353 2564 1369 2581
rect 1211 2547 1261 2564
rect 1061 2500 1261 2547
rect 1319 2547 1369 2564
rect 1469 2564 1485 2581
rect 1611 2581 1743 2597
rect 1611 2564 1627 2581
rect 1469 2547 1519 2564
rect 1319 2500 1519 2547
rect 1577 2547 1627 2564
rect 1727 2564 1743 2581
rect 1869 2581 2001 2597
rect 1869 2564 1885 2581
rect 1727 2547 1777 2564
rect 1577 2500 1777 2547
rect 1835 2547 1885 2564
rect 1985 2564 2001 2581
rect 2127 2581 2259 2597
rect 2127 2564 2143 2581
rect 1985 2547 2035 2564
rect 1835 2500 2035 2547
rect 2093 2547 2143 2564
rect 2243 2564 2259 2581
rect 2385 2581 2517 2597
rect 2385 2564 2401 2581
rect 2243 2547 2293 2564
rect 2093 2500 2293 2547
rect 2351 2547 2401 2564
rect 2501 2564 2517 2581
rect 2643 2581 2775 2597
rect 2643 2564 2659 2581
rect 2501 2547 2551 2564
rect 2351 2500 2551 2547
rect 2609 2547 2659 2564
rect 2759 2564 2775 2581
rect 2901 2581 3033 2597
rect 2901 2564 2917 2581
rect 2759 2547 2809 2564
rect 2609 2500 2809 2547
rect 2867 2547 2917 2564
rect 3017 2564 3033 2581
rect 3159 2581 3291 2597
rect 3159 2564 3175 2581
rect 3017 2547 3067 2564
rect 2867 2500 3067 2547
rect 3125 2547 3175 2564
rect 3275 2564 3291 2581
rect 3417 2581 3549 2597
rect 3417 2564 3433 2581
rect 3275 2547 3325 2564
rect 3125 2500 3325 2547
rect 3383 2547 3433 2564
rect 3533 2564 3549 2581
rect 3675 2581 3807 2597
rect 3675 2564 3691 2581
rect 3533 2547 3583 2564
rect 3383 2500 3583 2547
rect 3641 2547 3691 2564
rect 3791 2564 3807 2581
rect 3933 2581 4065 2597
rect 3933 2564 3949 2581
rect 3791 2547 3841 2564
rect 3641 2500 3841 2547
rect 3899 2547 3949 2564
rect 4049 2564 4065 2581
rect 4191 2581 4323 2597
rect 4191 2564 4207 2581
rect 4049 2547 4099 2564
rect 3899 2500 4099 2547
rect 4157 2547 4207 2564
rect 4307 2564 4323 2581
rect 4307 2547 4357 2564
rect 4157 2500 4357 2547
rect -4357 -2547 -4157 -2500
rect -4357 -2564 -4307 -2547
rect -4323 -2581 -4307 -2564
rect -4207 -2564 -4157 -2547
rect -4099 -2547 -3899 -2500
rect -4099 -2564 -4049 -2547
rect -4207 -2581 -4191 -2564
rect -4323 -2597 -4191 -2581
rect -4065 -2581 -4049 -2564
rect -3949 -2564 -3899 -2547
rect -3841 -2547 -3641 -2500
rect -3841 -2564 -3791 -2547
rect -3949 -2581 -3933 -2564
rect -4065 -2597 -3933 -2581
rect -3807 -2581 -3791 -2564
rect -3691 -2564 -3641 -2547
rect -3583 -2547 -3383 -2500
rect -3583 -2564 -3533 -2547
rect -3691 -2581 -3675 -2564
rect -3807 -2597 -3675 -2581
rect -3549 -2581 -3533 -2564
rect -3433 -2564 -3383 -2547
rect -3325 -2547 -3125 -2500
rect -3325 -2564 -3275 -2547
rect -3433 -2581 -3417 -2564
rect -3549 -2597 -3417 -2581
rect -3291 -2581 -3275 -2564
rect -3175 -2564 -3125 -2547
rect -3067 -2547 -2867 -2500
rect -3067 -2564 -3017 -2547
rect -3175 -2581 -3159 -2564
rect -3291 -2597 -3159 -2581
rect -3033 -2581 -3017 -2564
rect -2917 -2564 -2867 -2547
rect -2809 -2547 -2609 -2500
rect -2809 -2564 -2759 -2547
rect -2917 -2581 -2901 -2564
rect -3033 -2597 -2901 -2581
rect -2775 -2581 -2759 -2564
rect -2659 -2564 -2609 -2547
rect -2551 -2547 -2351 -2500
rect -2551 -2564 -2501 -2547
rect -2659 -2581 -2643 -2564
rect -2775 -2597 -2643 -2581
rect -2517 -2581 -2501 -2564
rect -2401 -2564 -2351 -2547
rect -2293 -2547 -2093 -2500
rect -2293 -2564 -2243 -2547
rect -2401 -2581 -2385 -2564
rect -2517 -2597 -2385 -2581
rect -2259 -2581 -2243 -2564
rect -2143 -2564 -2093 -2547
rect -2035 -2547 -1835 -2500
rect -2035 -2564 -1985 -2547
rect -2143 -2581 -2127 -2564
rect -2259 -2597 -2127 -2581
rect -2001 -2581 -1985 -2564
rect -1885 -2564 -1835 -2547
rect -1777 -2547 -1577 -2500
rect -1777 -2564 -1727 -2547
rect -1885 -2581 -1869 -2564
rect -2001 -2597 -1869 -2581
rect -1743 -2581 -1727 -2564
rect -1627 -2564 -1577 -2547
rect -1519 -2547 -1319 -2500
rect -1519 -2564 -1469 -2547
rect -1627 -2581 -1611 -2564
rect -1743 -2597 -1611 -2581
rect -1485 -2581 -1469 -2564
rect -1369 -2564 -1319 -2547
rect -1261 -2547 -1061 -2500
rect -1261 -2564 -1211 -2547
rect -1369 -2581 -1353 -2564
rect -1485 -2597 -1353 -2581
rect -1227 -2581 -1211 -2564
rect -1111 -2564 -1061 -2547
rect -1003 -2547 -803 -2500
rect -1003 -2564 -953 -2547
rect -1111 -2581 -1095 -2564
rect -1227 -2597 -1095 -2581
rect -969 -2581 -953 -2564
rect -853 -2564 -803 -2547
rect -745 -2547 -545 -2500
rect -745 -2564 -695 -2547
rect -853 -2581 -837 -2564
rect -969 -2597 -837 -2581
rect -711 -2581 -695 -2564
rect -595 -2564 -545 -2547
rect -487 -2547 -287 -2500
rect -487 -2564 -437 -2547
rect -595 -2581 -579 -2564
rect -711 -2597 -579 -2581
rect -453 -2581 -437 -2564
rect -337 -2564 -287 -2547
rect -229 -2547 -29 -2500
rect -229 -2564 -179 -2547
rect -337 -2581 -321 -2564
rect -453 -2597 -321 -2581
rect -195 -2581 -179 -2564
rect -79 -2564 -29 -2547
rect 29 -2547 229 -2500
rect 29 -2564 79 -2547
rect -79 -2581 -63 -2564
rect -195 -2597 -63 -2581
rect 63 -2581 79 -2564
rect 179 -2564 229 -2547
rect 287 -2547 487 -2500
rect 287 -2564 337 -2547
rect 179 -2581 195 -2564
rect 63 -2597 195 -2581
rect 321 -2581 337 -2564
rect 437 -2564 487 -2547
rect 545 -2547 745 -2500
rect 545 -2564 595 -2547
rect 437 -2581 453 -2564
rect 321 -2597 453 -2581
rect 579 -2581 595 -2564
rect 695 -2564 745 -2547
rect 803 -2547 1003 -2500
rect 803 -2564 853 -2547
rect 695 -2581 711 -2564
rect 579 -2597 711 -2581
rect 837 -2581 853 -2564
rect 953 -2564 1003 -2547
rect 1061 -2547 1261 -2500
rect 1061 -2564 1111 -2547
rect 953 -2581 969 -2564
rect 837 -2597 969 -2581
rect 1095 -2581 1111 -2564
rect 1211 -2564 1261 -2547
rect 1319 -2547 1519 -2500
rect 1319 -2564 1369 -2547
rect 1211 -2581 1227 -2564
rect 1095 -2597 1227 -2581
rect 1353 -2581 1369 -2564
rect 1469 -2564 1519 -2547
rect 1577 -2547 1777 -2500
rect 1577 -2564 1627 -2547
rect 1469 -2581 1485 -2564
rect 1353 -2597 1485 -2581
rect 1611 -2581 1627 -2564
rect 1727 -2564 1777 -2547
rect 1835 -2547 2035 -2500
rect 1835 -2564 1885 -2547
rect 1727 -2581 1743 -2564
rect 1611 -2597 1743 -2581
rect 1869 -2581 1885 -2564
rect 1985 -2564 2035 -2547
rect 2093 -2547 2293 -2500
rect 2093 -2564 2143 -2547
rect 1985 -2581 2001 -2564
rect 1869 -2597 2001 -2581
rect 2127 -2581 2143 -2564
rect 2243 -2564 2293 -2547
rect 2351 -2547 2551 -2500
rect 2351 -2564 2401 -2547
rect 2243 -2581 2259 -2564
rect 2127 -2597 2259 -2581
rect 2385 -2581 2401 -2564
rect 2501 -2564 2551 -2547
rect 2609 -2547 2809 -2500
rect 2609 -2564 2659 -2547
rect 2501 -2581 2517 -2564
rect 2385 -2597 2517 -2581
rect 2643 -2581 2659 -2564
rect 2759 -2564 2809 -2547
rect 2867 -2547 3067 -2500
rect 2867 -2564 2917 -2547
rect 2759 -2581 2775 -2564
rect 2643 -2597 2775 -2581
rect 2901 -2581 2917 -2564
rect 3017 -2564 3067 -2547
rect 3125 -2547 3325 -2500
rect 3125 -2564 3175 -2547
rect 3017 -2581 3033 -2564
rect 2901 -2597 3033 -2581
rect 3159 -2581 3175 -2564
rect 3275 -2564 3325 -2547
rect 3383 -2547 3583 -2500
rect 3383 -2564 3433 -2547
rect 3275 -2581 3291 -2564
rect 3159 -2597 3291 -2581
rect 3417 -2581 3433 -2564
rect 3533 -2564 3583 -2547
rect 3641 -2547 3841 -2500
rect 3641 -2564 3691 -2547
rect 3533 -2581 3549 -2564
rect 3417 -2597 3549 -2581
rect 3675 -2581 3691 -2564
rect 3791 -2564 3841 -2547
rect 3899 -2547 4099 -2500
rect 3899 -2564 3949 -2547
rect 3791 -2581 3807 -2564
rect 3675 -2597 3807 -2581
rect 3933 -2581 3949 -2564
rect 4049 -2564 4099 -2547
rect 4157 -2547 4357 -2500
rect 4157 -2564 4207 -2547
rect 4049 -2581 4065 -2564
rect 3933 -2597 4065 -2581
rect 4191 -2581 4207 -2564
rect 4307 -2564 4357 -2547
rect 4307 -2581 4323 -2564
rect 4191 -2597 4323 -2581
<< polycont >>
rect -4307 2547 -4207 2581
rect -4049 2547 -3949 2581
rect -3791 2547 -3691 2581
rect -3533 2547 -3433 2581
rect -3275 2547 -3175 2581
rect -3017 2547 -2917 2581
rect -2759 2547 -2659 2581
rect -2501 2547 -2401 2581
rect -2243 2547 -2143 2581
rect -1985 2547 -1885 2581
rect -1727 2547 -1627 2581
rect -1469 2547 -1369 2581
rect -1211 2547 -1111 2581
rect -953 2547 -853 2581
rect -695 2547 -595 2581
rect -437 2547 -337 2581
rect -179 2547 -79 2581
rect 79 2547 179 2581
rect 337 2547 437 2581
rect 595 2547 695 2581
rect 853 2547 953 2581
rect 1111 2547 1211 2581
rect 1369 2547 1469 2581
rect 1627 2547 1727 2581
rect 1885 2547 1985 2581
rect 2143 2547 2243 2581
rect 2401 2547 2501 2581
rect 2659 2547 2759 2581
rect 2917 2547 3017 2581
rect 3175 2547 3275 2581
rect 3433 2547 3533 2581
rect 3691 2547 3791 2581
rect 3949 2547 4049 2581
rect 4207 2547 4307 2581
rect -4307 -2581 -4207 -2547
rect -4049 -2581 -3949 -2547
rect -3791 -2581 -3691 -2547
rect -3533 -2581 -3433 -2547
rect -3275 -2581 -3175 -2547
rect -3017 -2581 -2917 -2547
rect -2759 -2581 -2659 -2547
rect -2501 -2581 -2401 -2547
rect -2243 -2581 -2143 -2547
rect -1985 -2581 -1885 -2547
rect -1727 -2581 -1627 -2547
rect -1469 -2581 -1369 -2547
rect -1211 -2581 -1111 -2547
rect -953 -2581 -853 -2547
rect -695 -2581 -595 -2547
rect -437 -2581 -337 -2547
rect -179 -2581 -79 -2547
rect 79 -2581 179 -2547
rect 337 -2581 437 -2547
rect 595 -2581 695 -2547
rect 853 -2581 953 -2547
rect 1111 -2581 1211 -2547
rect 1369 -2581 1469 -2547
rect 1627 -2581 1727 -2547
rect 1885 -2581 1985 -2547
rect 2143 -2581 2243 -2547
rect 2401 -2581 2501 -2547
rect 2659 -2581 2759 -2547
rect 2917 -2581 3017 -2547
rect 3175 -2581 3275 -2547
rect 3433 -2581 3533 -2547
rect 3691 -2581 3791 -2547
rect 3949 -2581 4049 -2547
rect 4207 -2581 4307 -2547
<< locali >>
rect -4537 2685 -4441 2719
rect 4441 2685 4537 2719
rect -4537 2623 -4503 2685
rect 4503 2623 4537 2685
rect -4323 2547 -4307 2581
rect -4207 2547 -4191 2581
rect -4065 2547 -4049 2581
rect -3949 2547 -3933 2581
rect -3807 2547 -3791 2581
rect -3691 2547 -3675 2581
rect -3549 2547 -3533 2581
rect -3433 2547 -3417 2581
rect -3291 2547 -3275 2581
rect -3175 2547 -3159 2581
rect -3033 2547 -3017 2581
rect -2917 2547 -2901 2581
rect -2775 2547 -2759 2581
rect -2659 2547 -2643 2581
rect -2517 2547 -2501 2581
rect -2401 2547 -2385 2581
rect -2259 2547 -2243 2581
rect -2143 2547 -2127 2581
rect -2001 2547 -1985 2581
rect -1885 2547 -1869 2581
rect -1743 2547 -1727 2581
rect -1627 2547 -1611 2581
rect -1485 2547 -1469 2581
rect -1369 2547 -1353 2581
rect -1227 2547 -1211 2581
rect -1111 2547 -1095 2581
rect -969 2547 -953 2581
rect -853 2547 -837 2581
rect -711 2547 -695 2581
rect -595 2547 -579 2581
rect -453 2547 -437 2581
rect -337 2547 -321 2581
rect -195 2547 -179 2581
rect -79 2547 -63 2581
rect 63 2547 79 2581
rect 179 2547 195 2581
rect 321 2547 337 2581
rect 437 2547 453 2581
rect 579 2547 595 2581
rect 695 2547 711 2581
rect 837 2547 853 2581
rect 953 2547 969 2581
rect 1095 2547 1111 2581
rect 1211 2547 1227 2581
rect 1353 2547 1369 2581
rect 1469 2547 1485 2581
rect 1611 2547 1627 2581
rect 1727 2547 1743 2581
rect 1869 2547 1885 2581
rect 1985 2547 2001 2581
rect 2127 2547 2143 2581
rect 2243 2547 2259 2581
rect 2385 2547 2401 2581
rect 2501 2547 2517 2581
rect 2643 2547 2659 2581
rect 2759 2547 2775 2581
rect 2901 2547 2917 2581
rect 3017 2547 3033 2581
rect 3159 2547 3175 2581
rect 3275 2547 3291 2581
rect 3417 2547 3433 2581
rect 3533 2547 3549 2581
rect 3675 2547 3691 2581
rect 3791 2547 3807 2581
rect 3933 2547 3949 2581
rect 4049 2547 4065 2581
rect 4191 2547 4207 2581
rect 4307 2547 4323 2581
rect -4403 2488 -4369 2504
rect -4403 -2504 -4369 -2488
rect -4145 2488 -4111 2504
rect -4145 -2504 -4111 -2488
rect -3887 2488 -3853 2504
rect -3887 -2504 -3853 -2488
rect -3629 2488 -3595 2504
rect -3629 -2504 -3595 -2488
rect -3371 2488 -3337 2504
rect -3371 -2504 -3337 -2488
rect -3113 2488 -3079 2504
rect -3113 -2504 -3079 -2488
rect -2855 2488 -2821 2504
rect -2855 -2504 -2821 -2488
rect -2597 2488 -2563 2504
rect -2597 -2504 -2563 -2488
rect -2339 2488 -2305 2504
rect -2339 -2504 -2305 -2488
rect -2081 2488 -2047 2504
rect -2081 -2504 -2047 -2488
rect -1823 2488 -1789 2504
rect -1823 -2504 -1789 -2488
rect -1565 2488 -1531 2504
rect -1565 -2504 -1531 -2488
rect -1307 2488 -1273 2504
rect -1307 -2504 -1273 -2488
rect -1049 2488 -1015 2504
rect -1049 -2504 -1015 -2488
rect -791 2488 -757 2504
rect -791 -2504 -757 -2488
rect -533 2488 -499 2504
rect -533 -2504 -499 -2488
rect -275 2488 -241 2504
rect -275 -2504 -241 -2488
rect -17 2488 17 2504
rect -17 -2504 17 -2488
rect 241 2488 275 2504
rect 241 -2504 275 -2488
rect 499 2488 533 2504
rect 499 -2504 533 -2488
rect 757 2488 791 2504
rect 757 -2504 791 -2488
rect 1015 2488 1049 2504
rect 1015 -2504 1049 -2488
rect 1273 2488 1307 2504
rect 1273 -2504 1307 -2488
rect 1531 2488 1565 2504
rect 1531 -2504 1565 -2488
rect 1789 2488 1823 2504
rect 1789 -2504 1823 -2488
rect 2047 2488 2081 2504
rect 2047 -2504 2081 -2488
rect 2305 2488 2339 2504
rect 2305 -2504 2339 -2488
rect 2563 2488 2597 2504
rect 2563 -2504 2597 -2488
rect 2821 2488 2855 2504
rect 2821 -2504 2855 -2488
rect 3079 2488 3113 2504
rect 3079 -2504 3113 -2488
rect 3337 2488 3371 2504
rect 3337 -2504 3371 -2488
rect 3595 2488 3629 2504
rect 3595 -2504 3629 -2488
rect 3853 2488 3887 2504
rect 3853 -2504 3887 -2488
rect 4111 2488 4145 2504
rect 4111 -2504 4145 -2488
rect 4369 2488 4403 2504
rect 4369 -2504 4403 -2488
rect -4323 -2581 -4307 -2547
rect -4207 -2581 -4191 -2547
rect -4065 -2581 -4049 -2547
rect -3949 -2581 -3933 -2547
rect -3807 -2581 -3791 -2547
rect -3691 -2581 -3675 -2547
rect -3549 -2581 -3533 -2547
rect -3433 -2581 -3417 -2547
rect -3291 -2581 -3275 -2547
rect -3175 -2581 -3159 -2547
rect -3033 -2581 -3017 -2547
rect -2917 -2581 -2901 -2547
rect -2775 -2581 -2759 -2547
rect -2659 -2581 -2643 -2547
rect -2517 -2581 -2501 -2547
rect -2401 -2581 -2385 -2547
rect -2259 -2581 -2243 -2547
rect -2143 -2581 -2127 -2547
rect -2001 -2581 -1985 -2547
rect -1885 -2581 -1869 -2547
rect -1743 -2581 -1727 -2547
rect -1627 -2581 -1611 -2547
rect -1485 -2581 -1469 -2547
rect -1369 -2581 -1353 -2547
rect -1227 -2581 -1211 -2547
rect -1111 -2581 -1095 -2547
rect -969 -2581 -953 -2547
rect -853 -2581 -837 -2547
rect -711 -2581 -695 -2547
rect -595 -2581 -579 -2547
rect -453 -2581 -437 -2547
rect -337 -2581 -321 -2547
rect -195 -2581 -179 -2547
rect -79 -2581 -63 -2547
rect 63 -2581 79 -2547
rect 179 -2581 195 -2547
rect 321 -2581 337 -2547
rect 437 -2581 453 -2547
rect 579 -2581 595 -2547
rect 695 -2581 711 -2547
rect 837 -2581 853 -2547
rect 953 -2581 969 -2547
rect 1095 -2581 1111 -2547
rect 1211 -2581 1227 -2547
rect 1353 -2581 1369 -2547
rect 1469 -2581 1485 -2547
rect 1611 -2581 1627 -2547
rect 1727 -2581 1743 -2547
rect 1869 -2581 1885 -2547
rect 1985 -2581 2001 -2547
rect 2127 -2581 2143 -2547
rect 2243 -2581 2259 -2547
rect 2385 -2581 2401 -2547
rect 2501 -2581 2517 -2547
rect 2643 -2581 2659 -2547
rect 2759 -2581 2775 -2547
rect 2901 -2581 2917 -2547
rect 3017 -2581 3033 -2547
rect 3159 -2581 3175 -2547
rect 3275 -2581 3291 -2547
rect 3417 -2581 3433 -2547
rect 3533 -2581 3549 -2547
rect 3675 -2581 3691 -2547
rect 3791 -2581 3807 -2547
rect 3933 -2581 3949 -2547
rect 4049 -2581 4065 -2547
rect 4191 -2581 4207 -2547
rect 4307 -2581 4323 -2547
rect -4537 -2685 -4503 -2623
rect 4503 -2685 4537 -2623
rect -4537 -2719 -4441 -2685
rect 4441 -2719 4537 -2685
<< viali >>
rect -4307 2547 -4207 2581
rect -4049 2547 -3949 2581
rect -3791 2547 -3691 2581
rect -3533 2547 -3433 2581
rect -3275 2547 -3175 2581
rect -3017 2547 -2917 2581
rect -2759 2547 -2659 2581
rect -2501 2547 -2401 2581
rect -2243 2547 -2143 2581
rect -1985 2547 -1885 2581
rect -1727 2547 -1627 2581
rect -1469 2547 -1369 2581
rect -1211 2547 -1111 2581
rect -953 2547 -853 2581
rect -695 2547 -595 2581
rect -437 2547 -337 2581
rect -179 2547 -79 2581
rect 79 2547 179 2581
rect 337 2547 437 2581
rect 595 2547 695 2581
rect 853 2547 953 2581
rect 1111 2547 1211 2581
rect 1369 2547 1469 2581
rect 1627 2547 1727 2581
rect 1885 2547 1985 2581
rect 2143 2547 2243 2581
rect 2401 2547 2501 2581
rect 2659 2547 2759 2581
rect 2917 2547 3017 2581
rect 3175 2547 3275 2581
rect 3433 2547 3533 2581
rect 3691 2547 3791 2581
rect 3949 2547 4049 2581
rect 4207 2547 4307 2581
rect -4403 -2488 -4369 2488
rect -4145 -2488 -4111 2488
rect -3887 -2488 -3853 2488
rect -3629 -2488 -3595 2488
rect -3371 -2488 -3337 2488
rect -3113 -2488 -3079 2488
rect -2855 -2488 -2821 2488
rect -2597 -2488 -2563 2488
rect -2339 -2488 -2305 2488
rect -2081 -2488 -2047 2488
rect -1823 -2488 -1789 2488
rect -1565 -2488 -1531 2488
rect -1307 -2488 -1273 2488
rect -1049 -2488 -1015 2488
rect -791 -2488 -757 2488
rect -533 -2488 -499 2488
rect -275 -2488 -241 2488
rect -17 -2488 17 2488
rect 241 -2488 275 2488
rect 499 -2488 533 2488
rect 757 -2488 791 2488
rect 1015 -2488 1049 2488
rect 1273 -2488 1307 2488
rect 1531 -2488 1565 2488
rect 1789 -2488 1823 2488
rect 2047 -2488 2081 2488
rect 2305 -2488 2339 2488
rect 2563 -2488 2597 2488
rect 2821 -2488 2855 2488
rect 3079 -2488 3113 2488
rect 3337 -2488 3371 2488
rect 3595 -2488 3629 2488
rect 3853 -2488 3887 2488
rect 4111 -2488 4145 2488
rect 4369 -2488 4403 2488
rect -4307 -2581 -4207 -2547
rect -4049 -2581 -3949 -2547
rect -3791 -2581 -3691 -2547
rect -3533 -2581 -3433 -2547
rect -3275 -2581 -3175 -2547
rect -3017 -2581 -2917 -2547
rect -2759 -2581 -2659 -2547
rect -2501 -2581 -2401 -2547
rect -2243 -2581 -2143 -2547
rect -1985 -2581 -1885 -2547
rect -1727 -2581 -1627 -2547
rect -1469 -2581 -1369 -2547
rect -1211 -2581 -1111 -2547
rect -953 -2581 -853 -2547
rect -695 -2581 -595 -2547
rect -437 -2581 -337 -2547
rect -179 -2581 -79 -2547
rect 79 -2581 179 -2547
rect 337 -2581 437 -2547
rect 595 -2581 695 -2547
rect 853 -2581 953 -2547
rect 1111 -2581 1211 -2547
rect 1369 -2581 1469 -2547
rect 1627 -2581 1727 -2547
rect 1885 -2581 1985 -2547
rect 2143 -2581 2243 -2547
rect 2401 -2581 2501 -2547
rect 2659 -2581 2759 -2547
rect 2917 -2581 3017 -2547
rect 3175 -2581 3275 -2547
rect 3433 -2581 3533 -2547
rect 3691 -2581 3791 -2547
rect 3949 -2581 4049 -2547
rect 4207 -2581 4307 -2547
<< metal1 >>
rect -4319 2581 -4195 2587
rect -4319 2547 -4307 2581
rect -4207 2547 -4195 2581
rect -4319 2541 -4195 2547
rect -4061 2581 -3937 2587
rect -4061 2547 -4049 2581
rect -3949 2547 -3937 2581
rect -4061 2541 -3937 2547
rect -3803 2581 -3679 2587
rect -3803 2547 -3791 2581
rect -3691 2547 -3679 2581
rect -3803 2541 -3679 2547
rect -3545 2581 -3421 2587
rect -3545 2547 -3533 2581
rect -3433 2547 -3421 2581
rect -3545 2541 -3421 2547
rect -3287 2581 -3163 2587
rect -3287 2547 -3275 2581
rect -3175 2547 -3163 2581
rect -3287 2541 -3163 2547
rect -3029 2581 -2905 2587
rect -3029 2547 -3017 2581
rect -2917 2547 -2905 2581
rect -3029 2541 -2905 2547
rect -2771 2581 -2647 2587
rect -2771 2547 -2759 2581
rect -2659 2547 -2647 2581
rect -2771 2541 -2647 2547
rect -2513 2581 -2389 2587
rect -2513 2547 -2501 2581
rect -2401 2547 -2389 2581
rect -2513 2541 -2389 2547
rect -2255 2581 -2131 2587
rect -2255 2547 -2243 2581
rect -2143 2547 -2131 2581
rect -2255 2541 -2131 2547
rect -1997 2581 -1873 2587
rect -1997 2547 -1985 2581
rect -1885 2547 -1873 2581
rect -1997 2541 -1873 2547
rect -1739 2581 -1615 2587
rect -1739 2547 -1727 2581
rect -1627 2547 -1615 2581
rect -1739 2541 -1615 2547
rect -1481 2581 -1357 2587
rect -1481 2547 -1469 2581
rect -1369 2547 -1357 2581
rect -1481 2541 -1357 2547
rect -1223 2581 -1099 2587
rect -1223 2547 -1211 2581
rect -1111 2547 -1099 2581
rect -1223 2541 -1099 2547
rect -965 2581 -841 2587
rect -965 2547 -953 2581
rect -853 2547 -841 2581
rect -965 2541 -841 2547
rect -707 2581 -583 2587
rect -707 2547 -695 2581
rect -595 2547 -583 2581
rect -707 2541 -583 2547
rect -449 2581 -325 2587
rect -449 2547 -437 2581
rect -337 2547 -325 2581
rect -449 2541 -325 2547
rect -191 2581 -67 2587
rect -191 2547 -179 2581
rect -79 2547 -67 2581
rect -191 2541 -67 2547
rect 67 2581 191 2587
rect 67 2547 79 2581
rect 179 2547 191 2581
rect 67 2541 191 2547
rect 325 2581 449 2587
rect 325 2547 337 2581
rect 437 2547 449 2581
rect 325 2541 449 2547
rect 583 2581 707 2587
rect 583 2547 595 2581
rect 695 2547 707 2581
rect 583 2541 707 2547
rect 841 2581 965 2587
rect 841 2547 853 2581
rect 953 2547 965 2581
rect 841 2541 965 2547
rect 1099 2581 1223 2587
rect 1099 2547 1111 2581
rect 1211 2547 1223 2581
rect 1099 2541 1223 2547
rect 1357 2581 1481 2587
rect 1357 2547 1369 2581
rect 1469 2547 1481 2581
rect 1357 2541 1481 2547
rect 1615 2581 1739 2587
rect 1615 2547 1627 2581
rect 1727 2547 1739 2581
rect 1615 2541 1739 2547
rect 1873 2581 1997 2587
rect 1873 2547 1885 2581
rect 1985 2547 1997 2581
rect 1873 2541 1997 2547
rect 2131 2581 2255 2587
rect 2131 2547 2143 2581
rect 2243 2547 2255 2581
rect 2131 2541 2255 2547
rect 2389 2581 2513 2587
rect 2389 2547 2401 2581
rect 2501 2547 2513 2581
rect 2389 2541 2513 2547
rect 2647 2581 2771 2587
rect 2647 2547 2659 2581
rect 2759 2547 2771 2581
rect 2647 2541 2771 2547
rect 2905 2581 3029 2587
rect 2905 2547 2917 2581
rect 3017 2547 3029 2581
rect 2905 2541 3029 2547
rect 3163 2581 3287 2587
rect 3163 2547 3175 2581
rect 3275 2547 3287 2581
rect 3163 2541 3287 2547
rect 3421 2581 3545 2587
rect 3421 2547 3433 2581
rect 3533 2547 3545 2581
rect 3421 2541 3545 2547
rect 3679 2581 3803 2587
rect 3679 2547 3691 2581
rect 3791 2547 3803 2581
rect 3679 2541 3803 2547
rect 3937 2581 4061 2587
rect 3937 2547 3949 2581
rect 4049 2547 4061 2581
rect 3937 2541 4061 2547
rect 4195 2581 4319 2587
rect 4195 2547 4207 2581
rect 4307 2547 4319 2581
rect 4195 2541 4319 2547
rect -4409 2488 -4363 2500
rect -4409 -2488 -4403 2488
rect -4369 -2488 -4363 2488
rect -4409 -2500 -4363 -2488
rect -4151 2488 -4105 2500
rect -4151 -2488 -4145 2488
rect -4111 -2488 -4105 2488
rect -4151 -2500 -4105 -2488
rect -3893 2488 -3847 2500
rect -3893 -2488 -3887 2488
rect -3853 -2488 -3847 2488
rect -3893 -2500 -3847 -2488
rect -3635 2488 -3589 2500
rect -3635 -2488 -3629 2488
rect -3595 -2488 -3589 2488
rect -3635 -2500 -3589 -2488
rect -3377 2488 -3331 2500
rect -3377 -2488 -3371 2488
rect -3337 -2488 -3331 2488
rect -3377 -2500 -3331 -2488
rect -3119 2488 -3073 2500
rect -3119 -2488 -3113 2488
rect -3079 -2488 -3073 2488
rect -3119 -2500 -3073 -2488
rect -2861 2488 -2815 2500
rect -2861 -2488 -2855 2488
rect -2821 -2488 -2815 2488
rect -2861 -2500 -2815 -2488
rect -2603 2488 -2557 2500
rect -2603 -2488 -2597 2488
rect -2563 -2488 -2557 2488
rect -2603 -2500 -2557 -2488
rect -2345 2488 -2299 2500
rect -2345 -2488 -2339 2488
rect -2305 -2488 -2299 2488
rect -2345 -2500 -2299 -2488
rect -2087 2488 -2041 2500
rect -2087 -2488 -2081 2488
rect -2047 -2488 -2041 2488
rect -2087 -2500 -2041 -2488
rect -1829 2488 -1783 2500
rect -1829 -2488 -1823 2488
rect -1789 -2488 -1783 2488
rect -1829 -2500 -1783 -2488
rect -1571 2488 -1525 2500
rect -1571 -2488 -1565 2488
rect -1531 -2488 -1525 2488
rect -1571 -2500 -1525 -2488
rect -1313 2488 -1267 2500
rect -1313 -2488 -1307 2488
rect -1273 -2488 -1267 2488
rect -1313 -2500 -1267 -2488
rect -1055 2488 -1009 2500
rect -1055 -2488 -1049 2488
rect -1015 -2488 -1009 2488
rect -1055 -2500 -1009 -2488
rect -797 2488 -751 2500
rect -797 -2488 -791 2488
rect -757 -2488 -751 2488
rect -797 -2500 -751 -2488
rect -539 2488 -493 2500
rect -539 -2488 -533 2488
rect -499 -2488 -493 2488
rect -539 -2500 -493 -2488
rect -281 2488 -235 2500
rect -281 -2488 -275 2488
rect -241 -2488 -235 2488
rect -281 -2500 -235 -2488
rect -23 2488 23 2500
rect -23 -2488 -17 2488
rect 17 -2488 23 2488
rect -23 -2500 23 -2488
rect 235 2488 281 2500
rect 235 -2488 241 2488
rect 275 -2488 281 2488
rect 235 -2500 281 -2488
rect 493 2488 539 2500
rect 493 -2488 499 2488
rect 533 -2488 539 2488
rect 493 -2500 539 -2488
rect 751 2488 797 2500
rect 751 -2488 757 2488
rect 791 -2488 797 2488
rect 751 -2500 797 -2488
rect 1009 2488 1055 2500
rect 1009 -2488 1015 2488
rect 1049 -2488 1055 2488
rect 1009 -2500 1055 -2488
rect 1267 2488 1313 2500
rect 1267 -2488 1273 2488
rect 1307 -2488 1313 2488
rect 1267 -2500 1313 -2488
rect 1525 2488 1571 2500
rect 1525 -2488 1531 2488
rect 1565 -2488 1571 2488
rect 1525 -2500 1571 -2488
rect 1783 2488 1829 2500
rect 1783 -2488 1789 2488
rect 1823 -2488 1829 2488
rect 1783 -2500 1829 -2488
rect 2041 2488 2087 2500
rect 2041 -2488 2047 2488
rect 2081 -2488 2087 2488
rect 2041 -2500 2087 -2488
rect 2299 2488 2345 2500
rect 2299 -2488 2305 2488
rect 2339 -2488 2345 2488
rect 2299 -2500 2345 -2488
rect 2557 2488 2603 2500
rect 2557 -2488 2563 2488
rect 2597 -2488 2603 2488
rect 2557 -2500 2603 -2488
rect 2815 2488 2861 2500
rect 2815 -2488 2821 2488
rect 2855 -2488 2861 2488
rect 2815 -2500 2861 -2488
rect 3073 2488 3119 2500
rect 3073 -2488 3079 2488
rect 3113 -2488 3119 2488
rect 3073 -2500 3119 -2488
rect 3331 2488 3377 2500
rect 3331 -2488 3337 2488
rect 3371 -2488 3377 2488
rect 3331 -2500 3377 -2488
rect 3589 2488 3635 2500
rect 3589 -2488 3595 2488
rect 3629 -2488 3635 2488
rect 3589 -2500 3635 -2488
rect 3847 2488 3893 2500
rect 3847 -2488 3853 2488
rect 3887 -2488 3893 2488
rect 3847 -2500 3893 -2488
rect 4105 2488 4151 2500
rect 4105 -2488 4111 2488
rect 4145 -2488 4151 2488
rect 4105 -2500 4151 -2488
rect 4363 2488 4409 2500
rect 4363 -2488 4369 2488
rect 4403 -2488 4409 2488
rect 4363 -2500 4409 -2488
rect -4319 -2547 -4195 -2541
rect -4319 -2581 -4307 -2547
rect -4207 -2581 -4195 -2547
rect -4319 -2587 -4195 -2581
rect -4061 -2547 -3937 -2541
rect -4061 -2581 -4049 -2547
rect -3949 -2581 -3937 -2547
rect -4061 -2587 -3937 -2581
rect -3803 -2547 -3679 -2541
rect -3803 -2581 -3791 -2547
rect -3691 -2581 -3679 -2547
rect -3803 -2587 -3679 -2581
rect -3545 -2547 -3421 -2541
rect -3545 -2581 -3533 -2547
rect -3433 -2581 -3421 -2547
rect -3545 -2587 -3421 -2581
rect -3287 -2547 -3163 -2541
rect -3287 -2581 -3275 -2547
rect -3175 -2581 -3163 -2547
rect -3287 -2587 -3163 -2581
rect -3029 -2547 -2905 -2541
rect -3029 -2581 -3017 -2547
rect -2917 -2581 -2905 -2547
rect -3029 -2587 -2905 -2581
rect -2771 -2547 -2647 -2541
rect -2771 -2581 -2759 -2547
rect -2659 -2581 -2647 -2547
rect -2771 -2587 -2647 -2581
rect -2513 -2547 -2389 -2541
rect -2513 -2581 -2501 -2547
rect -2401 -2581 -2389 -2547
rect -2513 -2587 -2389 -2581
rect -2255 -2547 -2131 -2541
rect -2255 -2581 -2243 -2547
rect -2143 -2581 -2131 -2547
rect -2255 -2587 -2131 -2581
rect -1997 -2547 -1873 -2541
rect -1997 -2581 -1985 -2547
rect -1885 -2581 -1873 -2547
rect -1997 -2587 -1873 -2581
rect -1739 -2547 -1615 -2541
rect -1739 -2581 -1727 -2547
rect -1627 -2581 -1615 -2547
rect -1739 -2587 -1615 -2581
rect -1481 -2547 -1357 -2541
rect -1481 -2581 -1469 -2547
rect -1369 -2581 -1357 -2547
rect -1481 -2587 -1357 -2581
rect -1223 -2547 -1099 -2541
rect -1223 -2581 -1211 -2547
rect -1111 -2581 -1099 -2547
rect -1223 -2587 -1099 -2581
rect -965 -2547 -841 -2541
rect -965 -2581 -953 -2547
rect -853 -2581 -841 -2547
rect -965 -2587 -841 -2581
rect -707 -2547 -583 -2541
rect -707 -2581 -695 -2547
rect -595 -2581 -583 -2547
rect -707 -2587 -583 -2581
rect -449 -2547 -325 -2541
rect -449 -2581 -437 -2547
rect -337 -2581 -325 -2547
rect -449 -2587 -325 -2581
rect -191 -2547 -67 -2541
rect -191 -2581 -179 -2547
rect -79 -2581 -67 -2547
rect -191 -2587 -67 -2581
rect 67 -2547 191 -2541
rect 67 -2581 79 -2547
rect 179 -2581 191 -2547
rect 67 -2587 191 -2581
rect 325 -2547 449 -2541
rect 325 -2581 337 -2547
rect 437 -2581 449 -2547
rect 325 -2587 449 -2581
rect 583 -2547 707 -2541
rect 583 -2581 595 -2547
rect 695 -2581 707 -2547
rect 583 -2587 707 -2581
rect 841 -2547 965 -2541
rect 841 -2581 853 -2547
rect 953 -2581 965 -2547
rect 841 -2587 965 -2581
rect 1099 -2547 1223 -2541
rect 1099 -2581 1111 -2547
rect 1211 -2581 1223 -2547
rect 1099 -2587 1223 -2581
rect 1357 -2547 1481 -2541
rect 1357 -2581 1369 -2547
rect 1469 -2581 1481 -2547
rect 1357 -2587 1481 -2581
rect 1615 -2547 1739 -2541
rect 1615 -2581 1627 -2547
rect 1727 -2581 1739 -2547
rect 1615 -2587 1739 -2581
rect 1873 -2547 1997 -2541
rect 1873 -2581 1885 -2547
rect 1985 -2581 1997 -2547
rect 1873 -2587 1997 -2581
rect 2131 -2547 2255 -2541
rect 2131 -2581 2143 -2547
rect 2243 -2581 2255 -2547
rect 2131 -2587 2255 -2581
rect 2389 -2547 2513 -2541
rect 2389 -2581 2401 -2547
rect 2501 -2581 2513 -2547
rect 2389 -2587 2513 -2581
rect 2647 -2547 2771 -2541
rect 2647 -2581 2659 -2547
rect 2759 -2581 2771 -2547
rect 2647 -2587 2771 -2581
rect 2905 -2547 3029 -2541
rect 2905 -2581 2917 -2547
rect 3017 -2581 3029 -2547
rect 2905 -2587 3029 -2581
rect 3163 -2547 3287 -2541
rect 3163 -2581 3175 -2547
rect 3275 -2581 3287 -2547
rect 3163 -2587 3287 -2581
rect 3421 -2547 3545 -2541
rect 3421 -2581 3433 -2547
rect 3533 -2581 3545 -2547
rect 3421 -2587 3545 -2581
rect 3679 -2547 3803 -2541
rect 3679 -2581 3691 -2547
rect 3791 -2581 3803 -2547
rect 3679 -2587 3803 -2581
rect 3937 -2547 4061 -2541
rect 3937 -2581 3949 -2547
rect 4049 -2581 4061 -2547
rect 3937 -2587 4061 -2581
rect 4195 -2547 4319 -2541
rect 4195 -2581 4207 -2547
rect 4307 -2581 4319 -2547
rect 4195 -2587 4319 -2581
<< properties >>
string FIXED_BBOX -4520 -2702 4520 2702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 25 l 1 m 1 nf 34 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

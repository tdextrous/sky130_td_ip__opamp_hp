magic
tech sky130A
magscale 1 2
timestamp 1713233716
<< nwell >>
rect -3583 -1615 3583 1615
<< mvpmos >>
rect -3325 118 -3125 1318
rect -3067 118 -2867 1318
rect -2809 118 -2609 1318
rect -2551 118 -2351 1318
rect -2293 118 -2093 1318
rect -2035 118 -1835 1318
rect -1777 118 -1577 1318
rect -1519 118 -1319 1318
rect -1261 118 -1061 1318
rect -1003 118 -803 1318
rect -745 118 -545 1318
rect -487 118 -287 1318
rect -229 118 -29 1318
rect 29 118 229 1318
rect 287 118 487 1318
rect 545 118 745 1318
rect 803 118 1003 1318
rect 1061 118 1261 1318
rect 1319 118 1519 1318
rect 1577 118 1777 1318
rect 1835 118 2035 1318
rect 2093 118 2293 1318
rect 2351 118 2551 1318
rect 2609 118 2809 1318
rect 2867 118 3067 1318
rect 3125 118 3325 1318
rect -3325 -1318 -3125 -118
rect -3067 -1318 -2867 -118
rect -2809 -1318 -2609 -118
rect -2551 -1318 -2351 -118
rect -2293 -1318 -2093 -118
rect -2035 -1318 -1835 -118
rect -1777 -1318 -1577 -118
rect -1519 -1318 -1319 -118
rect -1261 -1318 -1061 -118
rect -1003 -1318 -803 -118
rect -745 -1318 -545 -118
rect -487 -1318 -287 -118
rect -229 -1318 -29 -118
rect 29 -1318 229 -118
rect 287 -1318 487 -118
rect 545 -1318 745 -118
rect 803 -1318 1003 -118
rect 1061 -1318 1261 -118
rect 1319 -1318 1519 -118
rect 1577 -1318 1777 -118
rect 1835 -1318 2035 -118
rect 2093 -1318 2293 -118
rect 2351 -1318 2551 -118
rect 2609 -1318 2809 -118
rect 2867 -1318 3067 -118
rect 3125 -1318 3325 -118
<< mvpdiff >>
rect -3383 1306 -3325 1318
rect -3383 130 -3371 1306
rect -3337 130 -3325 1306
rect -3383 118 -3325 130
rect -3125 1306 -3067 1318
rect -3125 130 -3113 1306
rect -3079 130 -3067 1306
rect -3125 118 -3067 130
rect -2867 1306 -2809 1318
rect -2867 130 -2855 1306
rect -2821 130 -2809 1306
rect -2867 118 -2809 130
rect -2609 1306 -2551 1318
rect -2609 130 -2597 1306
rect -2563 130 -2551 1306
rect -2609 118 -2551 130
rect -2351 1306 -2293 1318
rect -2351 130 -2339 1306
rect -2305 130 -2293 1306
rect -2351 118 -2293 130
rect -2093 1306 -2035 1318
rect -2093 130 -2081 1306
rect -2047 130 -2035 1306
rect -2093 118 -2035 130
rect -1835 1306 -1777 1318
rect -1835 130 -1823 1306
rect -1789 130 -1777 1306
rect -1835 118 -1777 130
rect -1577 1306 -1519 1318
rect -1577 130 -1565 1306
rect -1531 130 -1519 1306
rect -1577 118 -1519 130
rect -1319 1306 -1261 1318
rect -1319 130 -1307 1306
rect -1273 130 -1261 1306
rect -1319 118 -1261 130
rect -1061 1306 -1003 1318
rect -1061 130 -1049 1306
rect -1015 130 -1003 1306
rect -1061 118 -1003 130
rect -803 1306 -745 1318
rect -803 130 -791 1306
rect -757 130 -745 1306
rect -803 118 -745 130
rect -545 1306 -487 1318
rect -545 130 -533 1306
rect -499 130 -487 1306
rect -545 118 -487 130
rect -287 1306 -229 1318
rect -287 130 -275 1306
rect -241 130 -229 1306
rect -287 118 -229 130
rect -29 1306 29 1318
rect -29 130 -17 1306
rect 17 130 29 1306
rect -29 118 29 130
rect 229 1306 287 1318
rect 229 130 241 1306
rect 275 130 287 1306
rect 229 118 287 130
rect 487 1306 545 1318
rect 487 130 499 1306
rect 533 130 545 1306
rect 487 118 545 130
rect 745 1306 803 1318
rect 745 130 757 1306
rect 791 130 803 1306
rect 745 118 803 130
rect 1003 1306 1061 1318
rect 1003 130 1015 1306
rect 1049 130 1061 1306
rect 1003 118 1061 130
rect 1261 1306 1319 1318
rect 1261 130 1273 1306
rect 1307 130 1319 1306
rect 1261 118 1319 130
rect 1519 1306 1577 1318
rect 1519 130 1531 1306
rect 1565 130 1577 1306
rect 1519 118 1577 130
rect 1777 1306 1835 1318
rect 1777 130 1789 1306
rect 1823 130 1835 1306
rect 1777 118 1835 130
rect 2035 1306 2093 1318
rect 2035 130 2047 1306
rect 2081 130 2093 1306
rect 2035 118 2093 130
rect 2293 1306 2351 1318
rect 2293 130 2305 1306
rect 2339 130 2351 1306
rect 2293 118 2351 130
rect 2551 1306 2609 1318
rect 2551 130 2563 1306
rect 2597 130 2609 1306
rect 2551 118 2609 130
rect 2809 1306 2867 1318
rect 2809 130 2821 1306
rect 2855 130 2867 1306
rect 2809 118 2867 130
rect 3067 1306 3125 1318
rect 3067 130 3079 1306
rect 3113 130 3125 1306
rect 3067 118 3125 130
rect 3325 1306 3383 1318
rect 3325 130 3337 1306
rect 3371 130 3383 1306
rect 3325 118 3383 130
rect -3383 -130 -3325 -118
rect -3383 -1306 -3371 -130
rect -3337 -1306 -3325 -130
rect -3383 -1318 -3325 -1306
rect -3125 -130 -3067 -118
rect -3125 -1306 -3113 -130
rect -3079 -1306 -3067 -130
rect -3125 -1318 -3067 -1306
rect -2867 -130 -2809 -118
rect -2867 -1306 -2855 -130
rect -2821 -1306 -2809 -130
rect -2867 -1318 -2809 -1306
rect -2609 -130 -2551 -118
rect -2609 -1306 -2597 -130
rect -2563 -1306 -2551 -130
rect -2609 -1318 -2551 -1306
rect -2351 -130 -2293 -118
rect -2351 -1306 -2339 -130
rect -2305 -1306 -2293 -130
rect -2351 -1318 -2293 -1306
rect -2093 -130 -2035 -118
rect -2093 -1306 -2081 -130
rect -2047 -1306 -2035 -130
rect -2093 -1318 -2035 -1306
rect -1835 -130 -1777 -118
rect -1835 -1306 -1823 -130
rect -1789 -1306 -1777 -130
rect -1835 -1318 -1777 -1306
rect -1577 -130 -1519 -118
rect -1577 -1306 -1565 -130
rect -1531 -1306 -1519 -130
rect -1577 -1318 -1519 -1306
rect -1319 -130 -1261 -118
rect -1319 -1306 -1307 -130
rect -1273 -1306 -1261 -130
rect -1319 -1318 -1261 -1306
rect -1061 -130 -1003 -118
rect -1061 -1306 -1049 -130
rect -1015 -1306 -1003 -130
rect -1061 -1318 -1003 -1306
rect -803 -130 -745 -118
rect -803 -1306 -791 -130
rect -757 -1306 -745 -130
rect -803 -1318 -745 -1306
rect -545 -130 -487 -118
rect -545 -1306 -533 -130
rect -499 -1306 -487 -130
rect -545 -1318 -487 -1306
rect -287 -130 -229 -118
rect -287 -1306 -275 -130
rect -241 -1306 -229 -130
rect -287 -1318 -229 -1306
rect -29 -130 29 -118
rect -29 -1306 -17 -130
rect 17 -1306 29 -130
rect -29 -1318 29 -1306
rect 229 -130 287 -118
rect 229 -1306 241 -130
rect 275 -1306 287 -130
rect 229 -1318 287 -1306
rect 487 -130 545 -118
rect 487 -1306 499 -130
rect 533 -1306 545 -130
rect 487 -1318 545 -1306
rect 745 -130 803 -118
rect 745 -1306 757 -130
rect 791 -1306 803 -130
rect 745 -1318 803 -1306
rect 1003 -130 1061 -118
rect 1003 -1306 1015 -130
rect 1049 -1306 1061 -130
rect 1003 -1318 1061 -1306
rect 1261 -130 1319 -118
rect 1261 -1306 1273 -130
rect 1307 -1306 1319 -130
rect 1261 -1318 1319 -1306
rect 1519 -130 1577 -118
rect 1519 -1306 1531 -130
rect 1565 -1306 1577 -130
rect 1519 -1318 1577 -1306
rect 1777 -130 1835 -118
rect 1777 -1306 1789 -130
rect 1823 -1306 1835 -130
rect 1777 -1318 1835 -1306
rect 2035 -130 2093 -118
rect 2035 -1306 2047 -130
rect 2081 -1306 2093 -130
rect 2035 -1318 2093 -1306
rect 2293 -130 2351 -118
rect 2293 -1306 2305 -130
rect 2339 -1306 2351 -130
rect 2293 -1318 2351 -1306
rect 2551 -130 2609 -118
rect 2551 -1306 2563 -130
rect 2597 -1306 2609 -130
rect 2551 -1318 2609 -1306
rect 2809 -130 2867 -118
rect 2809 -1306 2821 -130
rect 2855 -1306 2867 -130
rect 2809 -1318 2867 -1306
rect 3067 -130 3125 -118
rect 3067 -1306 3079 -130
rect 3113 -1306 3125 -130
rect 3067 -1318 3125 -1306
rect 3325 -130 3383 -118
rect 3325 -1306 3337 -130
rect 3371 -1306 3383 -130
rect 3325 -1318 3383 -1306
<< mvpdiffc >>
rect -3371 130 -3337 1306
rect -3113 130 -3079 1306
rect -2855 130 -2821 1306
rect -2597 130 -2563 1306
rect -2339 130 -2305 1306
rect -2081 130 -2047 1306
rect -1823 130 -1789 1306
rect -1565 130 -1531 1306
rect -1307 130 -1273 1306
rect -1049 130 -1015 1306
rect -791 130 -757 1306
rect -533 130 -499 1306
rect -275 130 -241 1306
rect -17 130 17 1306
rect 241 130 275 1306
rect 499 130 533 1306
rect 757 130 791 1306
rect 1015 130 1049 1306
rect 1273 130 1307 1306
rect 1531 130 1565 1306
rect 1789 130 1823 1306
rect 2047 130 2081 1306
rect 2305 130 2339 1306
rect 2563 130 2597 1306
rect 2821 130 2855 1306
rect 3079 130 3113 1306
rect 3337 130 3371 1306
rect -3371 -1306 -3337 -130
rect -3113 -1306 -3079 -130
rect -2855 -1306 -2821 -130
rect -2597 -1306 -2563 -130
rect -2339 -1306 -2305 -130
rect -2081 -1306 -2047 -130
rect -1823 -1306 -1789 -130
rect -1565 -1306 -1531 -130
rect -1307 -1306 -1273 -130
rect -1049 -1306 -1015 -130
rect -791 -1306 -757 -130
rect -533 -1306 -499 -130
rect -275 -1306 -241 -130
rect -17 -1306 17 -130
rect 241 -1306 275 -130
rect 499 -1306 533 -130
rect 757 -1306 791 -130
rect 1015 -1306 1049 -130
rect 1273 -1306 1307 -130
rect 1531 -1306 1565 -130
rect 1789 -1306 1823 -130
rect 2047 -1306 2081 -130
rect 2305 -1306 2339 -130
rect 2563 -1306 2597 -130
rect 2821 -1306 2855 -130
rect 3079 -1306 3113 -130
rect 3337 -1306 3371 -130
<< mvnsubdiff >>
rect -3517 1537 3517 1549
rect -3517 1503 -3409 1537
rect 3409 1503 3517 1537
rect -3517 1491 3517 1503
rect -3517 1441 -3459 1491
rect -3517 -1441 -3505 1441
rect -3471 -1441 -3459 1441
rect 3459 1441 3517 1491
rect -3517 -1491 -3459 -1441
rect 3459 -1441 3471 1441
rect 3505 -1441 3517 1441
rect 3459 -1491 3517 -1441
rect -3517 -1503 3517 -1491
rect -3517 -1537 -3409 -1503
rect 3409 -1537 3517 -1503
rect -3517 -1549 3517 -1537
<< mvnsubdiffcont >>
rect -3409 1503 3409 1537
rect -3505 -1441 -3471 1441
rect 3471 -1441 3505 1441
rect -3409 -1537 3409 -1503
<< poly >>
rect -3325 1399 -3125 1415
rect -3325 1365 -3309 1399
rect -3141 1365 -3125 1399
rect -3325 1318 -3125 1365
rect -3067 1399 -2867 1415
rect -3067 1365 -3051 1399
rect -2883 1365 -2867 1399
rect -3067 1318 -2867 1365
rect -2809 1399 -2609 1415
rect -2809 1365 -2793 1399
rect -2625 1365 -2609 1399
rect -2809 1318 -2609 1365
rect -2551 1399 -2351 1415
rect -2551 1365 -2535 1399
rect -2367 1365 -2351 1399
rect -2551 1318 -2351 1365
rect -2293 1399 -2093 1415
rect -2293 1365 -2277 1399
rect -2109 1365 -2093 1399
rect -2293 1318 -2093 1365
rect -2035 1399 -1835 1415
rect -2035 1365 -2019 1399
rect -1851 1365 -1835 1399
rect -2035 1318 -1835 1365
rect -1777 1399 -1577 1415
rect -1777 1365 -1761 1399
rect -1593 1365 -1577 1399
rect -1777 1318 -1577 1365
rect -1519 1399 -1319 1415
rect -1519 1365 -1503 1399
rect -1335 1365 -1319 1399
rect -1519 1318 -1319 1365
rect -1261 1399 -1061 1415
rect -1261 1365 -1245 1399
rect -1077 1365 -1061 1399
rect -1261 1318 -1061 1365
rect -1003 1399 -803 1415
rect -1003 1365 -987 1399
rect -819 1365 -803 1399
rect -1003 1318 -803 1365
rect -745 1399 -545 1415
rect -745 1365 -729 1399
rect -561 1365 -545 1399
rect -745 1318 -545 1365
rect -487 1399 -287 1415
rect -487 1365 -471 1399
rect -303 1365 -287 1399
rect -487 1318 -287 1365
rect -229 1399 -29 1415
rect -229 1365 -213 1399
rect -45 1365 -29 1399
rect -229 1318 -29 1365
rect 29 1399 229 1415
rect 29 1365 45 1399
rect 213 1365 229 1399
rect 29 1318 229 1365
rect 287 1399 487 1415
rect 287 1365 303 1399
rect 471 1365 487 1399
rect 287 1318 487 1365
rect 545 1399 745 1415
rect 545 1365 561 1399
rect 729 1365 745 1399
rect 545 1318 745 1365
rect 803 1399 1003 1415
rect 803 1365 819 1399
rect 987 1365 1003 1399
rect 803 1318 1003 1365
rect 1061 1399 1261 1415
rect 1061 1365 1077 1399
rect 1245 1365 1261 1399
rect 1061 1318 1261 1365
rect 1319 1399 1519 1415
rect 1319 1365 1335 1399
rect 1503 1365 1519 1399
rect 1319 1318 1519 1365
rect 1577 1399 1777 1415
rect 1577 1365 1593 1399
rect 1761 1365 1777 1399
rect 1577 1318 1777 1365
rect 1835 1399 2035 1415
rect 1835 1365 1851 1399
rect 2019 1365 2035 1399
rect 1835 1318 2035 1365
rect 2093 1399 2293 1415
rect 2093 1365 2109 1399
rect 2277 1365 2293 1399
rect 2093 1318 2293 1365
rect 2351 1399 2551 1415
rect 2351 1365 2367 1399
rect 2535 1365 2551 1399
rect 2351 1318 2551 1365
rect 2609 1399 2809 1415
rect 2609 1365 2625 1399
rect 2793 1365 2809 1399
rect 2609 1318 2809 1365
rect 2867 1399 3067 1415
rect 2867 1365 2883 1399
rect 3051 1365 3067 1399
rect 2867 1318 3067 1365
rect 3125 1399 3325 1415
rect 3125 1365 3141 1399
rect 3309 1365 3325 1399
rect 3125 1318 3325 1365
rect -3325 71 -3125 118
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3325 21 -3125 37
rect -3067 71 -2867 118
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -3067 21 -2867 37
rect -2809 71 -2609 118
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2809 21 -2609 37
rect -2551 71 -2351 118
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2551 21 -2351 37
rect -2293 71 -2093 118
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2293 21 -2093 37
rect -2035 71 -1835 118
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -2035 21 -1835 37
rect -1777 71 -1577 118
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1777 21 -1577 37
rect -1519 71 -1319 118
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1519 21 -1319 37
rect -1261 71 -1061 118
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1261 21 -1061 37
rect -1003 71 -803 118
rect -1003 37 -987 71
rect -819 37 -803 71
rect -1003 21 -803 37
rect -745 71 -545 118
rect -745 37 -729 71
rect -561 37 -545 71
rect -745 21 -545 37
rect -487 71 -287 118
rect -487 37 -471 71
rect -303 37 -287 71
rect -487 21 -287 37
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect 287 71 487 118
rect 287 37 303 71
rect 471 37 487 71
rect 287 21 487 37
rect 545 71 745 118
rect 545 37 561 71
rect 729 37 745 71
rect 545 21 745 37
rect 803 71 1003 118
rect 803 37 819 71
rect 987 37 1003 71
rect 803 21 1003 37
rect 1061 71 1261 118
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1061 21 1261 37
rect 1319 71 1519 118
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1319 21 1519 37
rect 1577 71 1777 118
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1577 21 1777 37
rect 1835 71 2035 118
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 1835 21 2035 37
rect 2093 71 2293 118
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2093 21 2293 37
rect 2351 71 2551 118
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2351 21 2551 37
rect 2609 71 2809 118
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2609 21 2809 37
rect 2867 71 3067 118
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 2867 21 3067 37
rect 3125 71 3325 118
rect 3125 37 3141 71
rect 3309 37 3325 71
rect 3125 21 3325 37
rect -3325 -37 -3125 -21
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3325 -118 -3125 -71
rect -3067 -37 -2867 -21
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -3067 -118 -2867 -71
rect -2809 -37 -2609 -21
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2809 -118 -2609 -71
rect -2551 -37 -2351 -21
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2551 -118 -2351 -71
rect -2293 -37 -2093 -21
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2293 -118 -2093 -71
rect -2035 -37 -1835 -21
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -2035 -118 -1835 -71
rect -1777 -37 -1577 -21
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1777 -118 -1577 -71
rect -1519 -37 -1319 -21
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1519 -118 -1319 -71
rect -1261 -37 -1061 -21
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1261 -118 -1061 -71
rect -1003 -37 -803 -21
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -1003 -118 -803 -71
rect -745 -37 -545 -21
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -745 -118 -545 -71
rect -487 -37 -287 -21
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -487 -118 -287 -71
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect 287 -37 487 -21
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 287 -118 487 -71
rect 545 -37 745 -21
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 545 -118 745 -71
rect 803 -37 1003 -21
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 803 -118 1003 -71
rect 1061 -37 1261 -21
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1061 -118 1261 -71
rect 1319 -37 1519 -21
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1319 -118 1519 -71
rect 1577 -37 1777 -21
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1577 -118 1777 -71
rect 1835 -37 2035 -21
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 1835 -118 2035 -71
rect 2093 -37 2293 -21
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2093 -118 2293 -71
rect 2351 -37 2551 -21
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2351 -118 2551 -71
rect 2609 -37 2809 -21
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2609 -118 2809 -71
rect 2867 -37 3067 -21
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 2867 -118 3067 -71
rect 3125 -37 3325 -21
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect 3125 -118 3325 -71
rect -3325 -1365 -3125 -1318
rect -3325 -1399 -3309 -1365
rect -3141 -1399 -3125 -1365
rect -3325 -1415 -3125 -1399
rect -3067 -1365 -2867 -1318
rect -3067 -1399 -3051 -1365
rect -2883 -1399 -2867 -1365
rect -3067 -1415 -2867 -1399
rect -2809 -1365 -2609 -1318
rect -2809 -1399 -2793 -1365
rect -2625 -1399 -2609 -1365
rect -2809 -1415 -2609 -1399
rect -2551 -1365 -2351 -1318
rect -2551 -1399 -2535 -1365
rect -2367 -1399 -2351 -1365
rect -2551 -1415 -2351 -1399
rect -2293 -1365 -2093 -1318
rect -2293 -1399 -2277 -1365
rect -2109 -1399 -2093 -1365
rect -2293 -1415 -2093 -1399
rect -2035 -1365 -1835 -1318
rect -2035 -1399 -2019 -1365
rect -1851 -1399 -1835 -1365
rect -2035 -1415 -1835 -1399
rect -1777 -1365 -1577 -1318
rect -1777 -1399 -1761 -1365
rect -1593 -1399 -1577 -1365
rect -1777 -1415 -1577 -1399
rect -1519 -1365 -1319 -1318
rect -1519 -1399 -1503 -1365
rect -1335 -1399 -1319 -1365
rect -1519 -1415 -1319 -1399
rect -1261 -1365 -1061 -1318
rect -1261 -1399 -1245 -1365
rect -1077 -1399 -1061 -1365
rect -1261 -1415 -1061 -1399
rect -1003 -1365 -803 -1318
rect -1003 -1399 -987 -1365
rect -819 -1399 -803 -1365
rect -1003 -1415 -803 -1399
rect -745 -1365 -545 -1318
rect -745 -1399 -729 -1365
rect -561 -1399 -545 -1365
rect -745 -1415 -545 -1399
rect -487 -1365 -287 -1318
rect -487 -1399 -471 -1365
rect -303 -1399 -287 -1365
rect -487 -1415 -287 -1399
rect -229 -1365 -29 -1318
rect -229 -1399 -213 -1365
rect -45 -1399 -29 -1365
rect -229 -1415 -29 -1399
rect 29 -1365 229 -1318
rect 29 -1399 45 -1365
rect 213 -1399 229 -1365
rect 29 -1415 229 -1399
rect 287 -1365 487 -1318
rect 287 -1399 303 -1365
rect 471 -1399 487 -1365
rect 287 -1415 487 -1399
rect 545 -1365 745 -1318
rect 545 -1399 561 -1365
rect 729 -1399 745 -1365
rect 545 -1415 745 -1399
rect 803 -1365 1003 -1318
rect 803 -1399 819 -1365
rect 987 -1399 1003 -1365
rect 803 -1415 1003 -1399
rect 1061 -1365 1261 -1318
rect 1061 -1399 1077 -1365
rect 1245 -1399 1261 -1365
rect 1061 -1415 1261 -1399
rect 1319 -1365 1519 -1318
rect 1319 -1399 1335 -1365
rect 1503 -1399 1519 -1365
rect 1319 -1415 1519 -1399
rect 1577 -1365 1777 -1318
rect 1577 -1399 1593 -1365
rect 1761 -1399 1777 -1365
rect 1577 -1415 1777 -1399
rect 1835 -1365 2035 -1318
rect 1835 -1399 1851 -1365
rect 2019 -1399 2035 -1365
rect 1835 -1415 2035 -1399
rect 2093 -1365 2293 -1318
rect 2093 -1399 2109 -1365
rect 2277 -1399 2293 -1365
rect 2093 -1415 2293 -1399
rect 2351 -1365 2551 -1318
rect 2351 -1399 2367 -1365
rect 2535 -1399 2551 -1365
rect 2351 -1415 2551 -1399
rect 2609 -1365 2809 -1318
rect 2609 -1399 2625 -1365
rect 2793 -1399 2809 -1365
rect 2609 -1415 2809 -1399
rect 2867 -1365 3067 -1318
rect 2867 -1399 2883 -1365
rect 3051 -1399 3067 -1365
rect 2867 -1415 3067 -1399
rect 3125 -1365 3325 -1318
rect 3125 -1399 3141 -1365
rect 3309 -1399 3325 -1365
rect 3125 -1415 3325 -1399
<< polycont >>
rect -3309 1365 -3141 1399
rect -3051 1365 -2883 1399
rect -2793 1365 -2625 1399
rect -2535 1365 -2367 1399
rect -2277 1365 -2109 1399
rect -2019 1365 -1851 1399
rect -1761 1365 -1593 1399
rect -1503 1365 -1335 1399
rect -1245 1365 -1077 1399
rect -987 1365 -819 1399
rect -729 1365 -561 1399
rect -471 1365 -303 1399
rect -213 1365 -45 1399
rect 45 1365 213 1399
rect 303 1365 471 1399
rect 561 1365 729 1399
rect 819 1365 987 1399
rect 1077 1365 1245 1399
rect 1335 1365 1503 1399
rect 1593 1365 1761 1399
rect 1851 1365 2019 1399
rect 2109 1365 2277 1399
rect 2367 1365 2535 1399
rect 2625 1365 2793 1399
rect 2883 1365 3051 1399
rect 3141 1365 3309 1399
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect -3309 -1399 -3141 -1365
rect -3051 -1399 -2883 -1365
rect -2793 -1399 -2625 -1365
rect -2535 -1399 -2367 -1365
rect -2277 -1399 -2109 -1365
rect -2019 -1399 -1851 -1365
rect -1761 -1399 -1593 -1365
rect -1503 -1399 -1335 -1365
rect -1245 -1399 -1077 -1365
rect -987 -1399 -819 -1365
rect -729 -1399 -561 -1365
rect -471 -1399 -303 -1365
rect -213 -1399 -45 -1365
rect 45 -1399 213 -1365
rect 303 -1399 471 -1365
rect 561 -1399 729 -1365
rect 819 -1399 987 -1365
rect 1077 -1399 1245 -1365
rect 1335 -1399 1503 -1365
rect 1593 -1399 1761 -1365
rect 1851 -1399 2019 -1365
rect 2109 -1399 2277 -1365
rect 2367 -1399 2535 -1365
rect 2625 -1399 2793 -1365
rect 2883 -1399 3051 -1365
rect 3141 -1399 3309 -1365
<< locali >>
rect -3505 1503 -3409 1537
rect 3409 1503 3505 1537
rect -3505 1441 -3471 1503
rect 3471 1441 3505 1503
rect -3325 1365 -3309 1399
rect -3141 1365 -3125 1399
rect -3067 1365 -3051 1399
rect -2883 1365 -2867 1399
rect -2809 1365 -2793 1399
rect -2625 1365 -2609 1399
rect -2551 1365 -2535 1399
rect -2367 1365 -2351 1399
rect -2293 1365 -2277 1399
rect -2109 1365 -2093 1399
rect -2035 1365 -2019 1399
rect -1851 1365 -1835 1399
rect -1777 1365 -1761 1399
rect -1593 1365 -1577 1399
rect -1519 1365 -1503 1399
rect -1335 1365 -1319 1399
rect -1261 1365 -1245 1399
rect -1077 1365 -1061 1399
rect -1003 1365 -987 1399
rect -819 1365 -803 1399
rect -745 1365 -729 1399
rect -561 1365 -545 1399
rect -487 1365 -471 1399
rect -303 1365 -287 1399
rect -229 1365 -213 1399
rect -45 1365 -29 1399
rect 29 1365 45 1399
rect 213 1365 229 1399
rect 287 1365 303 1399
rect 471 1365 487 1399
rect 545 1365 561 1399
rect 729 1365 745 1399
rect 803 1365 819 1399
rect 987 1365 1003 1399
rect 1061 1365 1077 1399
rect 1245 1365 1261 1399
rect 1319 1365 1335 1399
rect 1503 1365 1519 1399
rect 1577 1365 1593 1399
rect 1761 1365 1777 1399
rect 1835 1365 1851 1399
rect 2019 1365 2035 1399
rect 2093 1365 2109 1399
rect 2277 1365 2293 1399
rect 2351 1365 2367 1399
rect 2535 1365 2551 1399
rect 2609 1365 2625 1399
rect 2793 1365 2809 1399
rect 2867 1365 2883 1399
rect 3051 1365 3067 1399
rect 3125 1365 3141 1399
rect 3309 1365 3325 1399
rect -3371 1306 -3337 1322
rect -3371 114 -3337 130
rect -3113 1306 -3079 1322
rect -3113 114 -3079 130
rect -2855 1306 -2821 1322
rect -2855 114 -2821 130
rect -2597 1306 -2563 1322
rect -2597 114 -2563 130
rect -2339 1306 -2305 1322
rect -2339 114 -2305 130
rect -2081 1306 -2047 1322
rect -2081 114 -2047 130
rect -1823 1306 -1789 1322
rect -1823 114 -1789 130
rect -1565 1306 -1531 1322
rect -1565 114 -1531 130
rect -1307 1306 -1273 1322
rect -1307 114 -1273 130
rect -1049 1306 -1015 1322
rect -1049 114 -1015 130
rect -791 1306 -757 1322
rect -791 114 -757 130
rect -533 1306 -499 1322
rect -533 114 -499 130
rect -275 1306 -241 1322
rect -275 114 -241 130
rect -17 1306 17 1322
rect -17 114 17 130
rect 241 1306 275 1322
rect 241 114 275 130
rect 499 1306 533 1322
rect 499 114 533 130
rect 757 1306 791 1322
rect 757 114 791 130
rect 1015 1306 1049 1322
rect 1015 114 1049 130
rect 1273 1306 1307 1322
rect 1273 114 1307 130
rect 1531 1306 1565 1322
rect 1531 114 1565 130
rect 1789 1306 1823 1322
rect 1789 114 1823 130
rect 2047 1306 2081 1322
rect 2047 114 2081 130
rect 2305 1306 2339 1322
rect 2305 114 2339 130
rect 2563 1306 2597 1322
rect 2563 114 2597 130
rect 2821 1306 2855 1322
rect 2821 114 2855 130
rect 3079 1306 3113 1322
rect 3079 114 3113 130
rect 3337 1306 3371 1322
rect 3337 114 3371 130
rect -3325 37 -3309 71
rect -3141 37 -3125 71
rect -3067 37 -3051 71
rect -2883 37 -2867 71
rect -2809 37 -2793 71
rect -2625 37 -2609 71
rect -2551 37 -2535 71
rect -2367 37 -2351 71
rect -2293 37 -2277 71
rect -2109 37 -2093 71
rect -2035 37 -2019 71
rect -1851 37 -1835 71
rect -1777 37 -1761 71
rect -1593 37 -1577 71
rect -1519 37 -1503 71
rect -1335 37 -1319 71
rect -1261 37 -1245 71
rect -1077 37 -1061 71
rect -1003 37 -987 71
rect -819 37 -803 71
rect -745 37 -729 71
rect -561 37 -545 71
rect -487 37 -471 71
rect -303 37 -287 71
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect 287 37 303 71
rect 471 37 487 71
rect 545 37 561 71
rect 729 37 745 71
rect 803 37 819 71
rect 987 37 1003 71
rect 1061 37 1077 71
rect 1245 37 1261 71
rect 1319 37 1335 71
rect 1503 37 1519 71
rect 1577 37 1593 71
rect 1761 37 1777 71
rect 1835 37 1851 71
rect 2019 37 2035 71
rect 2093 37 2109 71
rect 2277 37 2293 71
rect 2351 37 2367 71
rect 2535 37 2551 71
rect 2609 37 2625 71
rect 2793 37 2809 71
rect 2867 37 2883 71
rect 3051 37 3067 71
rect 3125 37 3141 71
rect 3309 37 3325 71
rect -3325 -71 -3309 -37
rect -3141 -71 -3125 -37
rect -3067 -71 -3051 -37
rect -2883 -71 -2867 -37
rect -2809 -71 -2793 -37
rect -2625 -71 -2609 -37
rect -2551 -71 -2535 -37
rect -2367 -71 -2351 -37
rect -2293 -71 -2277 -37
rect -2109 -71 -2093 -37
rect -2035 -71 -2019 -37
rect -1851 -71 -1835 -37
rect -1777 -71 -1761 -37
rect -1593 -71 -1577 -37
rect -1519 -71 -1503 -37
rect -1335 -71 -1319 -37
rect -1261 -71 -1245 -37
rect -1077 -71 -1061 -37
rect -1003 -71 -987 -37
rect -819 -71 -803 -37
rect -745 -71 -729 -37
rect -561 -71 -545 -37
rect -487 -71 -471 -37
rect -303 -71 -287 -37
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 287 -71 303 -37
rect 471 -71 487 -37
rect 545 -71 561 -37
rect 729 -71 745 -37
rect 803 -71 819 -37
rect 987 -71 1003 -37
rect 1061 -71 1077 -37
rect 1245 -71 1261 -37
rect 1319 -71 1335 -37
rect 1503 -71 1519 -37
rect 1577 -71 1593 -37
rect 1761 -71 1777 -37
rect 1835 -71 1851 -37
rect 2019 -71 2035 -37
rect 2093 -71 2109 -37
rect 2277 -71 2293 -37
rect 2351 -71 2367 -37
rect 2535 -71 2551 -37
rect 2609 -71 2625 -37
rect 2793 -71 2809 -37
rect 2867 -71 2883 -37
rect 3051 -71 3067 -37
rect 3125 -71 3141 -37
rect 3309 -71 3325 -37
rect -3371 -130 -3337 -114
rect -3371 -1322 -3337 -1306
rect -3113 -130 -3079 -114
rect -3113 -1322 -3079 -1306
rect -2855 -130 -2821 -114
rect -2855 -1322 -2821 -1306
rect -2597 -130 -2563 -114
rect -2597 -1322 -2563 -1306
rect -2339 -130 -2305 -114
rect -2339 -1322 -2305 -1306
rect -2081 -130 -2047 -114
rect -2081 -1322 -2047 -1306
rect -1823 -130 -1789 -114
rect -1823 -1322 -1789 -1306
rect -1565 -130 -1531 -114
rect -1565 -1322 -1531 -1306
rect -1307 -130 -1273 -114
rect -1307 -1322 -1273 -1306
rect -1049 -130 -1015 -114
rect -1049 -1322 -1015 -1306
rect -791 -130 -757 -114
rect -791 -1322 -757 -1306
rect -533 -130 -499 -114
rect -533 -1322 -499 -1306
rect -275 -130 -241 -114
rect -275 -1322 -241 -1306
rect -17 -130 17 -114
rect -17 -1322 17 -1306
rect 241 -130 275 -114
rect 241 -1322 275 -1306
rect 499 -130 533 -114
rect 499 -1322 533 -1306
rect 757 -130 791 -114
rect 757 -1322 791 -1306
rect 1015 -130 1049 -114
rect 1015 -1322 1049 -1306
rect 1273 -130 1307 -114
rect 1273 -1322 1307 -1306
rect 1531 -130 1565 -114
rect 1531 -1322 1565 -1306
rect 1789 -130 1823 -114
rect 1789 -1322 1823 -1306
rect 2047 -130 2081 -114
rect 2047 -1322 2081 -1306
rect 2305 -130 2339 -114
rect 2305 -1322 2339 -1306
rect 2563 -130 2597 -114
rect 2563 -1322 2597 -1306
rect 2821 -130 2855 -114
rect 2821 -1322 2855 -1306
rect 3079 -130 3113 -114
rect 3079 -1322 3113 -1306
rect 3337 -130 3371 -114
rect 3337 -1322 3371 -1306
rect -3325 -1399 -3309 -1365
rect -3141 -1399 -3125 -1365
rect -3067 -1399 -3051 -1365
rect -2883 -1399 -2867 -1365
rect -2809 -1399 -2793 -1365
rect -2625 -1399 -2609 -1365
rect -2551 -1399 -2535 -1365
rect -2367 -1399 -2351 -1365
rect -2293 -1399 -2277 -1365
rect -2109 -1399 -2093 -1365
rect -2035 -1399 -2019 -1365
rect -1851 -1399 -1835 -1365
rect -1777 -1399 -1761 -1365
rect -1593 -1399 -1577 -1365
rect -1519 -1399 -1503 -1365
rect -1335 -1399 -1319 -1365
rect -1261 -1399 -1245 -1365
rect -1077 -1399 -1061 -1365
rect -1003 -1399 -987 -1365
rect -819 -1399 -803 -1365
rect -745 -1399 -729 -1365
rect -561 -1399 -545 -1365
rect -487 -1399 -471 -1365
rect -303 -1399 -287 -1365
rect -229 -1399 -213 -1365
rect -45 -1399 -29 -1365
rect 29 -1399 45 -1365
rect 213 -1399 229 -1365
rect 287 -1399 303 -1365
rect 471 -1399 487 -1365
rect 545 -1399 561 -1365
rect 729 -1399 745 -1365
rect 803 -1399 819 -1365
rect 987 -1399 1003 -1365
rect 1061 -1399 1077 -1365
rect 1245 -1399 1261 -1365
rect 1319 -1399 1335 -1365
rect 1503 -1399 1519 -1365
rect 1577 -1399 1593 -1365
rect 1761 -1399 1777 -1365
rect 1835 -1399 1851 -1365
rect 2019 -1399 2035 -1365
rect 2093 -1399 2109 -1365
rect 2277 -1399 2293 -1365
rect 2351 -1399 2367 -1365
rect 2535 -1399 2551 -1365
rect 2609 -1399 2625 -1365
rect 2793 -1399 2809 -1365
rect 2867 -1399 2883 -1365
rect 3051 -1399 3067 -1365
rect 3125 -1399 3141 -1365
rect 3309 -1399 3325 -1365
rect -3505 -1503 -3471 -1441
rect 3471 -1503 3505 -1441
rect -3505 -1537 -3409 -1503
rect 3409 -1537 3505 -1503
<< viali >>
rect -3309 1365 -3141 1399
rect -3051 1365 -2883 1399
rect -2793 1365 -2625 1399
rect -2535 1365 -2367 1399
rect -2277 1365 -2109 1399
rect -2019 1365 -1851 1399
rect -1761 1365 -1593 1399
rect -1503 1365 -1335 1399
rect -1245 1365 -1077 1399
rect -987 1365 -819 1399
rect -729 1365 -561 1399
rect -471 1365 -303 1399
rect -213 1365 -45 1399
rect 45 1365 213 1399
rect 303 1365 471 1399
rect 561 1365 729 1399
rect 819 1365 987 1399
rect 1077 1365 1245 1399
rect 1335 1365 1503 1399
rect 1593 1365 1761 1399
rect 1851 1365 2019 1399
rect 2109 1365 2277 1399
rect 2367 1365 2535 1399
rect 2625 1365 2793 1399
rect 2883 1365 3051 1399
rect 3141 1365 3309 1399
rect -3371 130 -3337 1306
rect -3113 130 -3079 1306
rect -2855 130 -2821 1306
rect -2597 130 -2563 1306
rect -2339 130 -2305 1306
rect -2081 130 -2047 1306
rect -1823 130 -1789 1306
rect -1565 130 -1531 1306
rect -1307 130 -1273 1306
rect -1049 130 -1015 1306
rect -791 130 -757 1306
rect -533 130 -499 1306
rect -275 130 -241 1306
rect -17 130 17 1306
rect 241 130 275 1306
rect 499 130 533 1306
rect 757 130 791 1306
rect 1015 130 1049 1306
rect 1273 130 1307 1306
rect 1531 130 1565 1306
rect 1789 130 1823 1306
rect 2047 130 2081 1306
rect 2305 130 2339 1306
rect 2563 130 2597 1306
rect 2821 130 2855 1306
rect 3079 130 3113 1306
rect 3337 130 3371 1306
rect -3309 37 -3141 71
rect -3051 37 -2883 71
rect -2793 37 -2625 71
rect -2535 37 -2367 71
rect -2277 37 -2109 71
rect -2019 37 -1851 71
rect -1761 37 -1593 71
rect -1503 37 -1335 71
rect -1245 37 -1077 71
rect -987 37 -819 71
rect -729 37 -561 71
rect -471 37 -303 71
rect -213 37 -45 71
rect 45 37 213 71
rect 303 37 471 71
rect 561 37 729 71
rect 819 37 987 71
rect 1077 37 1245 71
rect 1335 37 1503 71
rect 1593 37 1761 71
rect 1851 37 2019 71
rect 2109 37 2277 71
rect 2367 37 2535 71
rect 2625 37 2793 71
rect 2883 37 3051 71
rect 3141 37 3309 71
rect -3309 -71 -3141 -37
rect -3051 -71 -2883 -37
rect -2793 -71 -2625 -37
rect -2535 -71 -2367 -37
rect -2277 -71 -2109 -37
rect -2019 -71 -1851 -37
rect -1761 -71 -1593 -37
rect -1503 -71 -1335 -37
rect -1245 -71 -1077 -37
rect -987 -71 -819 -37
rect -729 -71 -561 -37
rect -471 -71 -303 -37
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect 303 -71 471 -37
rect 561 -71 729 -37
rect 819 -71 987 -37
rect 1077 -71 1245 -37
rect 1335 -71 1503 -37
rect 1593 -71 1761 -37
rect 1851 -71 2019 -37
rect 2109 -71 2277 -37
rect 2367 -71 2535 -37
rect 2625 -71 2793 -37
rect 2883 -71 3051 -37
rect 3141 -71 3309 -37
rect -3371 -1306 -3337 -130
rect -3113 -1306 -3079 -130
rect -2855 -1306 -2821 -130
rect -2597 -1306 -2563 -130
rect -2339 -1306 -2305 -130
rect -2081 -1306 -2047 -130
rect -1823 -1306 -1789 -130
rect -1565 -1306 -1531 -130
rect -1307 -1306 -1273 -130
rect -1049 -1306 -1015 -130
rect -791 -1306 -757 -130
rect -533 -1306 -499 -130
rect -275 -1306 -241 -130
rect -17 -1306 17 -130
rect 241 -1306 275 -130
rect 499 -1306 533 -130
rect 757 -1306 791 -130
rect 1015 -1306 1049 -130
rect 1273 -1306 1307 -130
rect 1531 -1306 1565 -130
rect 1789 -1306 1823 -130
rect 2047 -1306 2081 -130
rect 2305 -1306 2339 -130
rect 2563 -1306 2597 -130
rect 2821 -1306 2855 -130
rect 3079 -1306 3113 -130
rect 3337 -1306 3371 -130
rect -3309 -1399 -3141 -1365
rect -3051 -1399 -2883 -1365
rect -2793 -1399 -2625 -1365
rect -2535 -1399 -2367 -1365
rect -2277 -1399 -2109 -1365
rect -2019 -1399 -1851 -1365
rect -1761 -1399 -1593 -1365
rect -1503 -1399 -1335 -1365
rect -1245 -1399 -1077 -1365
rect -987 -1399 -819 -1365
rect -729 -1399 -561 -1365
rect -471 -1399 -303 -1365
rect -213 -1399 -45 -1365
rect 45 -1399 213 -1365
rect 303 -1399 471 -1365
rect 561 -1399 729 -1365
rect 819 -1399 987 -1365
rect 1077 -1399 1245 -1365
rect 1335 -1399 1503 -1365
rect 1593 -1399 1761 -1365
rect 1851 -1399 2019 -1365
rect 2109 -1399 2277 -1365
rect 2367 -1399 2535 -1365
rect 2625 -1399 2793 -1365
rect 2883 -1399 3051 -1365
rect 3141 -1399 3309 -1365
<< metal1 >>
rect -3321 1399 -3129 1405
rect -3321 1365 -3309 1399
rect -3141 1365 -3129 1399
rect -3321 1359 -3129 1365
rect -3063 1399 -2871 1405
rect -3063 1365 -3051 1399
rect -2883 1365 -2871 1399
rect -3063 1359 -2871 1365
rect -2805 1399 -2613 1405
rect -2805 1365 -2793 1399
rect -2625 1365 -2613 1399
rect -2805 1359 -2613 1365
rect -2547 1399 -2355 1405
rect -2547 1365 -2535 1399
rect -2367 1365 -2355 1399
rect -2547 1359 -2355 1365
rect -2289 1399 -2097 1405
rect -2289 1365 -2277 1399
rect -2109 1365 -2097 1399
rect -2289 1359 -2097 1365
rect -2031 1399 -1839 1405
rect -2031 1365 -2019 1399
rect -1851 1365 -1839 1399
rect -2031 1359 -1839 1365
rect -1773 1399 -1581 1405
rect -1773 1365 -1761 1399
rect -1593 1365 -1581 1399
rect -1773 1359 -1581 1365
rect -1515 1399 -1323 1405
rect -1515 1365 -1503 1399
rect -1335 1365 -1323 1399
rect -1515 1359 -1323 1365
rect -1257 1399 -1065 1405
rect -1257 1365 -1245 1399
rect -1077 1365 -1065 1399
rect -1257 1359 -1065 1365
rect -999 1399 -807 1405
rect -999 1365 -987 1399
rect -819 1365 -807 1399
rect -999 1359 -807 1365
rect -741 1399 -549 1405
rect -741 1365 -729 1399
rect -561 1365 -549 1399
rect -741 1359 -549 1365
rect -483 1399 -291 1405
rect -483 1365 -471 1399
rect -303 1365 -291 1399
rect -483 1359 -291 1365
rect -225 1399 -33 1405
rect -225 1365 -213 1399
rect -45 1365 -33 1399
rect -225 1359 -33 1365
rect 33 1399 225 1405
rect 33 1365 45 1399
rect 213 1365 225 1399
rect 33 1359 225 1365
rect 291 1399 483 1405
rect 291 1365 303 1399
rect 471 1365 483 1399
rect 291 1359 483 1365
rect 549 1399 741 1405
rect 549 1365 561 1399
rect 729 1365 741 1399
rect 549 1359 741 1365
rect 807 1399 999 1405
rect 807 1365 819 1399
rect 987 1365 999 1399
rect 807 1359 999 1365
rect 1065 1399 1257 1405
rect 1065 1365 1077 1399
rect 1245 1365 1257 1399
rect 1065 1359 1257 1365
rect 1323 1399 1515 1405
rect 1323 1365 1335 1399
rect 1503 1365 1515 1399
rect 1323 1359 1515 1365
rect 1581 1399 1773 1405
rect 1581 1365 1593 1399
rect 1761 1365 1773 1399
rect 1581 1359 1773 1365
rect 1839 1399 2031 1405
rect 1839 1365 1851 1399
rect 2019 1365 2031 1399
rect 1839 1359 2031 1365
rect 2097 1399 2289 1405
rect 2097 1365 2109 1399
rect 2277 1365 2289 1399
rect 2097 1359 2289 1365
rect 2355 1399 2547 1405
rect 2355 1365 2367 1399
rect 2535 1365 2547 1399
rect 2355 1359 2547 1365
rect 2613 1399 2805 1405
rect 2613 1365 2625 1399
rect 2793 1365 2805 1399
rect 2613 1359 2805 1365
rect 2871 1399 3063 1405
rect 2871 1365 2883 1399
rect 3051 1365 3063 1399
rect 2871 1359 3063 1365
rect 3129 1399 3321 1405
rect 3129 1365 3141 1399
rect 3309 1365 3321 1399
rect 3129 1359 3321 1365
rect -3377 1306 -3331 1318
rect -3377 130 -3371 1306
rect -3337 130 -3331 1306
rect -3377 118 -3331 130
rect -3119 1306 -3073 1318
rect -3119 130 -3113 1306
rect -3079 130 -3073 1306
rect -3119 118 -3073 130
rect -2861 1306 -2815 1318
rect -2861 130 -2855 1306
rect -2821 130 -2815 1306
rect -2861 118 -2815 130
rect -2603 1306 -2557 1318
rect -2603 130 -2597 1306
rect -2563 130 -2557 1306
rect -2603 118 -2557 130
rect -2345 1306 -2299 1318
rect -2345 130 -2339 1306
rect -2305 130 -2299 1306
rect -2345 118 -2299 130
rect -2087 1306 -2041 1318
rect -2087 130 -2081 1306
rect -2047 130 -2041 1306
rect -2087 118 -2041 130
rect -1829 1306 -1783 1318
rect -1829 130 -1823 1306
rect -1789 130 -1783 1306
rect -1829 118 -1783 130
rect -1571 1306 -1525 1318
rect -1571 130 -1565 1306
rect -1531 130 -1525 1306
rect -1571 118 -1525 130
rect -1313 1306 -1267 1318
rect -1313 130 -1307 1306
rect -1273 130 -1267 1306
rect -1313 118 -1267 130
rect -1055 1306 -1009 1318
rect -1055 130 -1049 1306
rect -1015 130 -1009 1306
rect -1055 118 -1009 130
rect -797 1306 -751 1318
rect -797 130 -791 1306
rect -757 130 -751 1306
rect -797 118 -751 130
rect -539 1306 -493 1318
rect -539 130 -533 1306
rect -499 130 -493 1306
rect -539 118 -493 130
rect -281 1306 -235 1318
rect -281 130 -275 1306
rect -241 130 -235 1306
rect -281 118 -235 130
rect -23 1306 23 1318
rect -23 130 -17 1306
rect 17 130 23 1306
rect -23 118 23 130
rect 235 1306 281 1318
rect 235 130 241 1306
rect 275 130 281 1306
rect 235 118 281 130
rect 493 1306 539 1318
rect 493 130 499 1306
rect 533 130 539 1306
rect 493 118 539 130
rect 751 1306 797 1318
rect 751 130 757 1306
rect 791 130 797 1306
rect 751 118 797 130
rect 1009 1306 1055 1318
rect 1009 130 1015 1306
rect 1049 130 1055 1306
rect 1009 118 1055 130
rect 1267 1306 1313 1318
rect 1267 130 1273 1306
rect 1307 130 1313 1306
rect 1267 118 1313 130
rect 1525 1306 1571 1318
rect 1525 130 1531 1306
rect 1565 130 1571 1306
rect 1525 118 1571 130
rect 1783 1306 1829 1318
rect 1783 130 1789 1306
rect 1823 130 1829 1306
rect 1783 118 1829 130
rect 2041 1306 2087 1318
rect 2041 130 2047 1306
rect 2081 130 2087 1306
rect 2041 118 2087 130
rect 2299 1306 2345 1318
rect 2299 130 2305 1306
rect 2339 130 2345 1306
rect 2299 118 2345 130
rect 2557 1306 2603 1318
rect 2557 130 2563 1306
rect 2597 130 2603 1306
rect 2557 118 2603 130
rect 2815 1306 2861 1318
rect 2815 130 2821 1306
rect 2855 130 2861 1306
rect 2815 118 2861 130
rect 3073 1306 3119 1318
rect 3073 130 3079 1306
rect 3113 130 3119 1306
rect 3073 118 3119 130
rect 3331 1306 3377 1318
rect 3331 130 3337 1306
rect 3371 130 3377 1306
rect 3331 118 3377 130
rect -3321 71 -3129 77
rect -3321 37 -3309 71
rect -3141 37 -3129 71
rect -3321 31 -3129 37
rect -3063 71 -2871 77
rect -3063 37 -3051 71
rect -2883 37 -2871 71
rect -3063 31 -2871 37
rect -2805 71 -2613 77
rect -2805 37 -2793 71
rect -2625 37 -2613 71
rect -2805 31 -2613 37
rect -2547 71 -2355 77
rect -2547 37 -2535 71
rect -2367 37 -2355 71
rect -2547 31 -2355 37
rect -2289 71 -2097 77
rect -2289 37 -2277 71
rect -2109 37 -2097 71
rect -2289 31 -2097 37
rect -2031 71 -1839 77
rect -2031 37 -2019 71
rect -1851 37 -1839 71
rect -2031 31 -1839 37
rect -1773 71 -1581 77
rect -1773 37 -1761 71
rect -1593 37 -1581 71
rect -1773 31 -1581 37
rect -1515 71 -1323 77
rect -1515 37 -1503 71
rect -1335 37 -1323 71
rect -1515 31 -1323 37
rect -1257 71 -1065 77
rect -1257 37 -1245 71
rect -1077 37 -1065 71
rect -1257 31 -1065 37
rect -999 71 -807 77
rect -999 37 -987 71
rect -819 37 -807 71
rect -999 31 -807 37
rect -741 71 -549 77
rect -741 37 -729 71
rect -561 37 -549 71
rect -741 31 -549 37
rect -483 71 -291 77
rect -483 37 -471 71
rect -303 37 -291 71
rect -483 31 -291 37
rect -225 71 -33 77
rect -225 37 -213 71
rect -45 37 -33 71
rect -225 31 -33 37
rect 33 71 225 77
rect 33 37 45 71
rect 213 37 225 71
rect 33 31 225 37
rect 291 71 483 77
rect 291 37 303 71
rect 471 37 483 71
rect 291 31 483 37
rect 549 71 741 77
rect 549 37 561 71
rect 729 37 741 71
rect 549 31 741 37
rect 807 71 999 77
rect 807 37 819 71
rect 987 37 999 71
rect 807 31 999 37
rect 1065 71 1257 77
rect 1065 37 1077 71
rect 1245 37 1257 71
rect 1065 31 1257 37
rect 1323 71 1515 77
rect 1323 37 1335 71
rect 1503 37 1515 71
rect 1323 31 1515 37
rect 1581 71 1773 77
rect 1581 37 1593 71
rect 1761 37 1773 71
rect 1581 31 1773 37
rect 1839 71 2031 77
rect 1839 37 1851 71
rect 2019 37 2031 71
rect 1839 31 2031 37
rect 2097 71 2289 77
rect 2097 37 2109 71
rect 2277 37 2289 71
rect 2097 31 2289 37
rect 2355 71 2547 77
rect 2355 37 2367 71
rect 2535 37 2547 71
rect 2355 31 2547 37
rect 2613 71 2805 77
rect 2613 37 2625 71
rect 2793 37 2805 71
rect 2613 31 2805 37
rect 2871 71 3063 77
rect 2871 37 2883 71
rect 3051 37 3063 71
rect 2871 31 3063 37
rect 3129 71 3321 77
rect 3129 37 3141 71
rect 3309 37 3321 71
rect 3129 31 3321 37
rect -3321 -37 -3129 -31
rect -3321 -71 -3309 -37
rect -3141 -71 -3129 -37
rect -3321 -77 -3129 -71
rect -3063 -37 -2871 -31
rect -3063 -71 -3051 -37
rect -2883 -71 -2871 -37
rect -3063 -77 -2871 -71
rect -2805 -37 -2613 -31
rect -2805 -71 -2793 -37
rect -2625 -71 -2613 -37
rect -2805 -77 -2613 -71
rect -2547 -37 -2355 -31
rect -2547 -71 -2535 -37
rect -2367 -71 -2355 -37
rect -2547 -77 -2355 -71
rect -2289 -37 -2097 -31
rect -2289 -71 -2277 -37
rect -2109 -71 -2097 -37
rect -2289 -77 -2097 -71
rect -2031 -37 -1839 -31
rect -2031 -71 -2019 -37
rect -1851 -71 -1839 -37
rect -2031 -77 -1839 -71
rect -1773 -37 -1581 -31
rect -1773 -71 -1761 -37
rect -1593 -71 -1581 -37
rect -1773 -77 -1581 -71
rect -1515 -37 -1323 -31
rect -1515 -71 -1503 -37
rect -1335 -71 -1323 -37
rect -1515 -77 -1323 -71
rect -1257 -37 -1065 -31
rect -1257 -71 -1245 -37
rect -1077 -71 -1065 -37
rect -1257 -77 -1065 -71
rect -999 -37 -807 -31
rect -999 -71 -987 -37
rect -819 -71 -807 -37
rect -999 -77 -807 -71
rect -741 -37 -549 -31
rect -741 -71 -729 -37
rect -561 -71 -549 -37
rect -741 -77 -549 -71
rect -483 -37 -291 -31
rect -483 -71 -471 -37
rect -303 -71 -291 -37
rect -483 -77 -291 -71
rect -225 -37 -33 -31
rect -225 -71 -213 -37
rect -45 -71 -33 -37
rect -225 -77 -33 -71
rect 33 -37 225 -31
rect 33 -71 45 -37
rect 213 -71 225 -37
rect 33 -77 225 -71
rect 291 -37 483 -31
rect 291 -71 303 -37
rect 471 -71 483 -37
rect 291 -77 483 -71
rect 549 -37 741 -31
rect 549 -71 561 -37
rect 729 -71 741 -37
rect 549 -77 741 -71
rect 807 -37 999 -31
rect 807 -71 819 -37
rect 987 -71 999 -37
rect 807 -77 999 -71
rect 1065 -37 1257 -31
rect 1065 -71 1077 -37
rect 1245 -71 1257 -37
rect 1065 -77 1257 -71
rect 1323 -37 1515 -31
rect 1323 -71 1335 -37
rect 1503 -71 1515 -37
rect 1323 -77 1515 -71
rect 1581 -37 1773 -31
rect 1581 -71 1593 -37
rect 1761 -71 1773 -37
rect 1581 -77 1773 -71
rect 1839 -37 2031 -31
rect 1839 -71 1851 -37
rect 2019 -71 2031 -37
rect 1839 -77 2031 -71
rect 2097 -37 2289 -31
rect 2097 -71 2109 -37
rect 2277 -71 2289 -37
rect 2097 -77 2289 -71
rect 2355 -37 2547 -31
rect 2355 -71 2367 -37
rect 2535 -71 2547 -37
rect 2355 -77 2547 -71
rect 2613 -37 2805 -31
rect 2613 -71 2625 -37
rect 2793 -71 2805 -37
rect 2613 -77 2805 -71
rect 2871 -37 3063 -31
rect 2871 -71 2883 -37
rect 3051 -71 3063 -37
rect 2871 -77 3063 -71
rect 3129 -37 3321 -31
rect 3129 -71 3141 -37
rect 3309 -71 3321 -37
rect 3129 -77 3321 -71
rect -3377 -130 -3331 -118
rect -3377 -1306 -3371 -130
rect -3337 -1306 -3331 -130
rect -3377 -1318 -3331 -1306
rect -3119 -130 -3073 -118
rect -3119 -1306 -3113 -130
rect -3079 -1306 -3073 -130
rect -3119 -1318 -3073 -1306
rect -2861 -130 -2815 -118
rect -2861 -1306 -2855 -130
rect -2821 -1306 -2815 -130
rect -2861 -1318 -2815 -1306
rect -2603 -130 -2557 -118
rect -2603 -1306 -2597 -130
rect -2563 -1306 -2557 -130
rect -2603 -1318 -2557 -1306
rect -2345 -130 -2299 -118
rect -2345 -1306 -2339 -130
rect -2305 -1306 -2299 -130
rect -2345 -1318 -2299 -1306
rect -2087 -130 -2041 -118
rect -2087 -1306 -2081 -130
rect -2047 -1306 -2041 -130
rect -2087 -1318 -2041 -1306
rect -1829 -130 -1783 -118
rect -1829 -1306 -1823 -130
rect -1789 -1306 -1783 -130
rect -1829 -1318 -1783 -1306
rect -1571 -130 -1525 -118
rect -1571 -1306 -1565 -130
rect -1531 -1306 -1525 -130
rect -1571 -1318 -1525 -1306
rect -1313 -130 -1267 -118
rect -1313 -1306 -1307 -130
rect -1273 -1306 -1267 -130
rect -1313 -1318 -1267 -1306
rect -1055 -130 -1009 -118
rect -1055 -1306 -1049 -130
rect -1015 -1306 -1009 -130
rect -1055 -1318 -1009 -1306
rect -797 -130 -751 -118
rect -797 -1306 -791 -130
rect -757 -1306 -751 -130
rect -797 -1318 -751 -1306
rect -539 -130 -493 -118
rect -539 -1306 -533 -130
rect -499 -1306 -493 -130
rect -539 -1318 -493 -1306
rect -281 -130 -235 -118
rect -281 -1306 -275 -130
rect -241 -1306 -235 -130
rect -281 -1318 -235 -1306
rect -23 -130 23 -118
rect -23 -1306 -17 -130
rect 17 -1306 23 -130
rect -23 -1318 23 -1306
rect 235 -130 281 -118
rect 235 -1306 241 -130
rect 275 -1306 281 -130
rect 235 -1318 281 -1306
rect 493 -130 539 -118
rect 493 -1306 499 -130
rect 533 -1306 539 -130
rect 493 -1318 539 -1306
rect 751 -130 797 -118
rect 751 -1306 757 -130
rect 791 -1306 797 -130
rect 751 -1318 797 -1306
rect 1009 -130 1055 -118
rect 1009 -1306 1015 -130
rect 1049 -1306 1055 -130
rect 1009 -1318 1055 -1306
rect 1267 -130 1313 -118
rect 1267 -1306 1273 -130
rect 1307 -1306 1313 -130
rect 1267 -1318 1313 -1306
rect 1525 -130 1571 -118
rect 1525 -1306 1531 -130
rect 1565 -1306 1571 -130
rect 1525 -1318 1571 -1306
rect 1783 -130 1829 -118
rect 1783 -1306 1789 -130
rect 1823 -1306 1829 -130
rect 1783 -1318 1829 -1306
rect 2041 -130 2087 -118
rect 2041 -1306 2047 -130
rect 2081 -1306 2087 -130
rect 2041 -1318 2087 -1306
rect 2299 -130 2345 -118
rect 2299 -1306 2305 -130
rect 2339 -1306 2345 -130
rect 2299 -1318 2345 -1306
rect 2557 -130 2603 -118
rect 2557 -1306 2563 -130
rect 2597 -1306 2603 -130
rect 2557 -1318 2603 -1306
rect 2815 -130 2861 -118
rect 2815 -1306 2821 -130
rect 2855 -1306 2861 -130
rect 2815 -1318 2861 -1306
rect 3073 -130 3119 -118
rect 3073 -1306 3079 -130
rect 3113 -1306 3119 -130
rect 3073 -1318 3119 -1306
rect 3331 -130 3377 -118
rect 3331 -1306 3337 -130
rect 3371 -1306 3377 -130
rect 3331 -1318 3377 -1306
rect -3321 -1365 -3129 -1359
rect -3321 -1399 -3309 -1365
rect -3141 -1399 -3129 -1365
rect -3321 -1405 -3129 -1399
rect -3063 -1365 -2871 -1359
rect -3063 -1399 -3051 -1365
rect -2883 -1399 -2871 -1365
rect -3063 -1405 -2871 -1399
rect -2805 -1365 -2613 -1359
rect -2805 -1399 -2793 -1365
rect -2625 -1399 -2613 -1365
rect -2805 -1405 -2613 -1399
rect -2547 -1365 -2355 -1359
rect -2547 -1399 -2535 -1365
rect -2367 -1399 -2355 -1365
rect -2547 -1405 -2355 -1399
rect -2289 -1365 -2097 -1359
rect -2289 -1399 -2277 -1365
rect -2109 -1399 -2097 -1365
rect -2289 -1405 -2097 -1399
rect -2031 -1365 -1839 -1359
rect -2031 -1399 -2019 -1365
rect -1851 -1399 -1839 -1365
rect -2031 -1405 -1839 -1399
rect -1773 -1365 -1581 -1359
rect -1773 -1399 -1761 -1365
rect -1593 -1399 -1581 -1365
rect -1773 -1405 -1581 -1399
rect -1515 -1365 -1323 -1359
rect -1515 -1399 -1503 -1365
rect -1335 -1399 -1323 -1365
rect -1515 -1405 -1323 -1399
rect -1257 -1365 -1065 -1359
rect -1257 -1399 -1245 -1365
rect -1077 -1399 -1065 -1365
rect -1257 -1405 -1065 -1399
rect -999 -1365 -807 -1359
rect -999 -1399 -987 -1365
rect -819 -1399 -807 -1365
rect -999 -1405 -807 -1399
rect -741 -1365 -549 -1359
rect -741 -1399 -729 -1365
rect -561 -1399 -549 -1365
rect -741 -1405 -549 -1399
rect -483 -1365 -291 -1359
rect -483 -1399 -471 -1365
rect -303 -1399 -291 -1365
rect -483 -1405 -291 -1399
rect -225 -1365 -33 -1359
rect -225 -1399 -213 -1365
rect -45 -1399 -33 -1365
rect -225 -1405 -33 -1399
rect 33 -1365 225 -1359
rect 33 -1399 45 -1365
rect 213 -1399 225 -1365
rect 33 -1405 225 -1399
rect 291 -1365 483 -1359
rect 291 -1399 303 -1365
rect 471 -1399 483 -1365
rect 291 -1405 483 -1399
rect 549 -1365 741 -1359
rect 549 -1399 561 -1365
rect 729 -1399 741 -1365
rect 549 -1405 741 -1399
rect 807 -1365 999 -1359
rect 807 -1399 819 -1365
rect 987 -1399 999 -1365
rect 807 -1405 999 -1399
rect 1065 -1365 1257 -1359
rect 1065 -1399 1077 -1365
rect 1245 -1399 1257 -1365
rect 1065 -1405 1257 -1399
rect 1323 -1365 1515 -1359
rect 1323 -1399 1335 -1365
rect 1503 -1399 1515 -1365
rect 1323 -1405 1515 -1399
rect 1581 -1365 1773 -1359
rect 1581 -1399 1593 -1365
rect 1761 -1399 1773 -1365
rect 1581 -1405 1773 -1399
rect 1839 -1365 2031 -1359
rect 1839 -1399 1851 -1365
rect 2019 -1399 2031 -1365
rect 1839 -1405 2031 -1399
rect 2097 -1365 2289 -1359
rect 2097 -1399 2109 -1365
rect 2277 -1399 2289 -1365
rect 2097 -1405 2289 -1399
rect 2355 -1365 2547 -1359
rect 2355 -1399 2367 -1365
rect 2535 -1399 2547 -1365
rect 2355 -1405 2547 -1399
rect 2613 -1365 2805 -1359
rect 2613 -1399 2625 -1365
rect 2793 -1399 2805 -1365
rect 2613 -1405 2805 -1399
rect 2871 -1365 3063 -1359
rect 2871 -1399 2883 -1365
rect 3051 -1399 3063 -1365
rect 2871 -1405 3063 -1399
rect 3129 -1365 3321 -1359
rect 3129 -1399 3141 -1365
rect 3309 -1399 3321 -1365
rect 3129 -1405 3321 -1399
<< properties >>
string FIXED_BBOX -3488 -1520 3488 1520
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6 l 1 m 2 nf 26 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

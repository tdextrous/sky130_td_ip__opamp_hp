magic
tech sky130A
magscale 1 2
timestamp 1713297702
<< pwell >>
rect -4069 -708 4069 708
<< mvnmos >>
rect -3841 -450 -3641 450
rect -3583 -450 -3383 450
rect -3325 -450 -3125 450
rect -3067 -450 -2867 450
rect -2809 -450 -2609 450
rect -2551 -450 -2351 450
rect -2293 -450 -2093 450
rect -2035 -450 -1835 450
rect -1777 -450 -1577 450
rect -1519 -450 -1319 450
rect -1261 -450 -1061 450
rect -1003 -450 -803 450
rect -745 -450 -545 450
rect -487 -450 -287 450
rect -229 -450 -29 450
rect 29 -450 229 450
rect 287 -450 487 450
rect 545 -450 745 450
rect 803 -450 1003 450
rect 1061 -450 1261 450
rect 1319 -450 1519 450
rect 1577 -450 1777 450
rect 1835 -450 2035 450
rect 2093 -450 2293 450
rect 2351 -450 2551 450
rect 2609 -450 2809 450
rect 2867 -450 3067 450
rect 3125 -450 3325 450
rect 3383 -450 3583 450
rect 3641 -450 3841 450
<< mvndiff >>
rect -3899 438 -3841 450
rect -3899 -438 -3887 438
rect -3853 -438 -3841 438
rect -3899 -450 -3841 -438
rect -3641 438 -3583 450
rect -3641 -438 -3629 438
rect -3595 -438 -3583 438
rect -3641 -450 -3583 -438
rect -3383 438 -3325 450
rect -3383 -438 -3371 438
rect -3337 -438 -3325 438
rect -3383 -450 -3325 -438
rect -3125 438 -3067 450
rect -3125 -438 -3113 438
rect -3079 -438 -3067 438
rect -3125 -450 -3067 -438
rect -2867 438 -2809 450
rect -2867 -438 -2855 438
rect -2821 -438 -2809 438
rect -2867 -450 -2809 -438
rect -2609 438 -2551 450
rect -2609 -438 -2597 438
rect -2563 -438 -2551 438
rect -2609 -450 -2551 -438
rect -2351 438 -2293 450
rect -2351 -438 -2339 438
rect -2305 -438 -2293 438
rect -2351 -450 -2293 -438
rect -2093 438 -2035 450
rect -2093 -438 -2081 438
rect -2047 -438 -2035 438
rect -2093 -450 -2035 -438
rect -1835 438 -1777 450
rect -1835 -438 -1823 438
rect -1789 -438 -1777 438
rect -1835 -450 -1777 -438
rect -1577 438 -1519 450
rect -1577 -438 -1565 438
rect -1531 -438 -1519 438
rect -1577 -450 -1519 -438
rect -1319 438 -1261 450
rect -1319 -438 -1307 438
rect -1273 -438 -1261 438
rect -1319 -450 -1261 -438
rect -1061 438 -1003 450
rect -1061 -438 -1049 438
rect -1015 -438 -1003 438
rect -1061 -450 -1003 -438
rect -803 438 -745 450
rect -803 -438 -791 438
rect -757 -438 -745 438
rect -803 -450 -745 -438
rect -545 438 -487 450
rect -545 -438 -533 438
rect -499 -438 -487 438
rect -545 -450 -487 -438
rect -287 438 -229 450
rect -287 -438 -275 438
rect -241 -438 -229 438
rect -287 -450 -229 -438
rect -29 438 29 450
rect -29 -438 -17 438
rect 17 -438 29 438
rect -29 -450 29 -438
rect 229 438 287 450
rect 229 -438 241 438
rect 275 -438 287 438
rect 229 -450 287 -438
rect 487 438 545 450
rect 487 -438 499 438
rect 533 -438 545 438
rect 487 -450 545 -438
rect 745 438 803 450
rect 745 -438 757 438
rect 791 -438 803 438
rect 745 -450 803 -438
rect 1003 438 1061 450
rect 1003 -438 1015 438
rect 1049 -438 1061 438
rect 1003 -450 1061 -438
rect 1261 438 1319 450
rect 1261 -438 1273 438
rect 1307 -438 1319 438
rect 1261 -450 1319 -438
rect 1519 438 1577 450
rect 1519 -438 1531 438
rect 1565 -438 1577 438
rect 1519 -450 1577 -438
rect 1777 438 1835 450
rect 1777 -438 1789 438
rect 1823 -438 1835 438
rect 1777 -450 1835 -438
rect 2035 438 2093 450
rect 2035 -438 2047 438
rect 2081 -438 2093 438
rect 2035 -450 2093 -438
rect 2293 438 2351 450
rect 2293 -438 2305 438
rect 2339 -438 2351 438
rect 2293 -450 2351 -438
rect 2551 438 2609 450
rect 2551 -438 2563 438
rect 2597 -438 2609 438
rect 2551 -450 2609 -438
rect 2809 438 2867 450
rect 2809 -438 2821 438
rect 2855 -438 2867 438
rect 2809 -450 2867 -438
rect 3067 438 3125 450
rect 3067 -438 3079 438
rect 3113 -438 3125 438
rect 3067 -450 3125 -438
rect 3325 438 3383 450
rect 3325 -438 3337 438
rect 3371 -438 3383 438
rect 3325 -450 3383 -438
rect 3583 438 3641 450
rect 3583 -438 3595 438
rect 3629 -438 3641 438
rect 3583 -450 3641 -438
rect 3841 438 3899 450
rect 3841 -438 3853 438
rect 3887 -438 3899 438
rect 3841 -450 3899 -438
<< mvndiffc >>
rect -3887 -438 -3853 438
rect -3629 -438 -3595 438
rect -3371 -438 -3337 438
rect -3113 -438 -3079 438
rect -2855 -438 -2821 438
rect -2597 -438 -2563 438
rect -2339 -438 -2305 438
rect -2081 -438 -2047 438
rect -1823 -438 -1789 438
rect -1565 -438 -1531 438
rect -1307 -438 -1273 438
rect -1049 -438 -1015 438
rect -791 -438 -757 438
rect -533 -438 -499 438
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
rect 499 -438 533 438
rect 757 -438 791 438
rect 1015 -438 1049 438
rect 1273 -438 1307 438
rect 1531 -438 1565 438
rect 1789 -438 1823 438
rect 2047 -438 2081 438
rect 2305 -438 2339 438
rect 2563 -438 2597 438
rect 2821 -438 2855 438
rect 3079 -438 3113 438
rect 3337 -438 3371 438
rect 3595 -438 3629 438
rect 3853 -438 3887 438
<< mvpsubdiff >>
rect -4033 660 4033 672
rect -4033 626 -3925 660
rect 3925 626 4033 660
rect -4033 614 4033 626
rect -4033 564 -3975 614
rect -4033 -564 -4021 564
rect -3987 -564 -3975 564
rect 3975 564 4033 614
rect -4033 -614 -3975 -564
rect 3975 -564 3987 564
rect 4021 -564 4033 564
rect 3975 -614 4033 -564
rect -4033 -626 4033 -614
rect -4033 -660 -3925 -626
rect 3925 -660 4033 -626
rect -4033 -672 4033 -660
<< mvpsubdiffcont >>
rect -3925 626 3925 660
rect -4021 -564 -3987 564
rect 3987 -564 4021 564
rect -3925 -660 3925 -626
<< poly >>
rect -3807 522 -3675 538
rect -3807 505 -3791 522
rect -3841 488 -3791 505
rect -3691 505 -3675 522
rect -3549 522 -3417 538
rect -3549 505 -3533 522
rect -3691 488 -3641 505
rect -3841 450 -3641 488
rect -3583 488 -3533 505
rect -3433 505 -3417 522
rect -3291 522 -3159 538
rect -3291 505 -3275 522
rect -3433 488 -3383 505
rect -3583 450 -3383 488
rect -3325 488 -3275 505
rect -3175 505 -3159 522
rect -3033 522 -2901 538
rect -3033 505 -3017 522
rect -3175 488 -3125 505
rect -3325 450 -3125 488
rect -3067 488 -3017 505
rect -2917 505 -2901 522
rect -2775 522 -2643 538
rect -2775 505 -2759 522
rect -2917 488 -2867 505
rect -3067 450 -2867 488
rect -2809 488 -2759 505
rect -2659 505 -2643 522
rect -2517 522 -2385 538
rect -2517 505 -2501 522
rect -2659 488 -2609 505
rect -2809 450 -2609 488
rect -2551 488 -2501 505
rect -2401 505 -2385 522
rect -2259 522 -2127 538
rect -2259 505 -2243 522
rect -2401 488 -2351 505
rect -2551 450 -2351 488
rect -2293 488 -2243 505
rect -2143 505 -2127 522
rect -2001 522 -1869 538
rect -2001 505 -1985 522
rect -2143 488 -2093 505
rect -2293 450 -2093 488
rect -2035 488 -1985 505
rect -1885 505 -1869 522
rect -1743 522 -1611 538
rect -1743 505 -1727 522
rect -1885 488 -1835 505
rect -2035 450 -1835 488
rect -1777 488 -1727 505
rect -1627 505 -1611 522
rect -1485 522 -1353 538
rect -1485 505 -1469 522
rect -1627 488 -1577 505
rect -1777 450 -1577 488
rect -1519 488 -1469 505
rect -1369 505 -1353 522
rect -1227 522 -1095 538
rect -1227 505 -1211 522
rect -1369 488 -1319 505
rect -1519 450 -1319 488
rect -1261 488 -1211 505
rect -1111 505 -1095 522
rect -969 522 -837 538
rect -969 505 -953 522
rect -1111 488 -1061 505
rect -1261 450 -1061 488
rect -1003 488 -953 505
rect -853 505 -837 522
rect -711 522 -579 538
rect -711 505 -695 522
rect -853 488 -803 505
rect -1003 450 -803 488
rect -745 488 -695 505
rect -595 505 -579 522
rect -453 522 -321 538
rect -453 505 -437 522
rect -595 488 -545 505
rect -745 450 -545 488
rect -487 488 -437 505
rect -337 505 -321 522
rect -195 522 -63 538
rect -195 505 -179 522
rect -337 488 -287 505
rect -487 450 -287 488
rect -229 488 -179 505
rect -79 505 -63 522
rect 63 522 195 538
rect 63 505 79 522
rect -79 488 -29 505
rect -229 450 -29 488
rect 29 488 79 505
rect 179 505 195 522
rect 321 522 453 538
rect 321 505 337 522
rect 179 488 229 505
rect 29 450 229 488
rect 287 488 337 505
rect 437 505 453 522
rect 579 522 711 538
rect 579 505 595 522
rect 437 488 487 505
rect 287 450 487 488
rect 545 488 595 505
rect 695 505 711 522
rect 837 522 969 538
rect 837 505 853 522
rect 695 488 745 505
rect 545 450 745 488
rect 803 488 853 505
rect 953 505 969 522
rect 1095 522 1227 538
rect 1095 505 1111 522
rect 953 488 1003 505
rect 803 450 1003 488
rect 1061 488 1111 505
rect 1211 505 1227 522
rect 1353 522 1485 538
rect 1353 505 1369 522
rect 1211 488 1261 505
rect 1061 450 1261 488
rect 1319 488 1369 505
rect 1469 505 1485 522
rect 1611 522 1743 538
rect 1611 505 1627 522
rect 1469 488 1519 505
rect 1319 450 1519 488
rect 1577 488 1627 505
rect 1727 505 1743 522
rect 1869 522 2001 538
rect 1869 505 1885 522
rect 1727 488 1777 505
rect 1577 450 1777 488
rect 1835 488 1885 505
rect 1985 505 2001 522
rect 2127 522 2259 538
rect 2127 505 2143 522
rect 1985 488 2035 505
rect 1835 450 2035 488
rect 2093 488 2143 505
rect 2243 505 2259 522
rect 2385 522 2517 538
rect 2385 505 2401 522
rect 2243 488 2293 505
rect 2093 450 2293 488
rect 2351 488 2401 505
rect 2501 505 2517 522
rect 2643 522 2775 538
rect 2643 505 2659 522
rect 2501 488 2551 505
rect 2351 450 2551 488
rect 2609 488 2659 505
rect 2759 505 2775 522
rect 2901 522 3033 538
rect 2901 505 2917 522
rect 2759 488 2809 505
rect 2609 450 2809 488
rect 2867 488 2917 505
rect 3017 505 3033 522
rect 3159 522 3291 538
rect 3159 505 3175 522
rect 3017 488 3067 505
rect 2867 450 3067 488
rect 3125 488 3175 505
rect 3275 505 3291 522
rect 3417 522 3549 538
rect 3417 505 3433 522
rect 3275 488 3325 505
rect 3125 450 3325 488
rect 3383 488 3433 505
rect 3533 505 3549 522
rect 3675 522 3807 538
rect 3675 505 3691 522
rect 3533 488 3583 505
rect 3383 450 3583 488
rect 3641 488 3691 505
rect 3791 505 3807 522
rect 3791 488 3841 505
rect 3641 450 3841 488
rect -3841 -488 -3641 -450
rect -3841 -505 -3791 -488
rect -3807 -522 -3791 -505
rect -3691 -505 -3641 -488
rect -3583 -488 -3383 -450
rect -3583 -505 -3533 -488
rect -3691 -522 -3675 -505
rect -3807 -538 -3675 -522
rect -3549 -522 -3533 -505
rect -3433 -505 -3383 -488
rect -3325 -488 -3125 -450
rect -3325 -505 -3275 -488
rect -3433 -522 -3417 -505
rect -3549 -538 -3417 -522
rect -3291 -522 -3275 -505
rect -3175 -505 -3125 -488
rect -3067 -488 -2867 -450
rect -3067 -505 -3017 -488
rect -3175 -522 -3159 -505
rect -3291 -538 -3159 -522
rect -3033 -522 -3017 -505
rect -2917 -505 -2867 -488
rect -2809 -488 -2609 -450
rect -2809 -505 -2759 -488
rect -2917 -522 -2901 -505
rect -3033 -538 -2901 -522
rect -2775 -522 -2759 -505
rect -2659 -505 -2609 -488
rect -2551 -488 -2351 -450
rect -2551 -505 -2501 -488
rect -2659 -522 -2643 -505
rect -2775 -538 -2643 -522
rect -2517 -522 -2501 -505
rect -2401 -505 -2351 -488
rect -2293 -488 -2093 -450
rect -2293 -505 -2243 -488
rect -2401 -522 -2385 -505
rect -2517 -538 -2385 -522
rect -2259 -522 -2243 -505
rect -2143 -505 -2093 -488
rect -2035 -488 -1835 -450
rect -2035 -505 -1985 -488
rect -2143 -522 -2127 -505
rect -2259 -538 -2127 -522
rect -2001 -522 -1985 -505
rect -1885 -505 -1835 -488
rect -1777 -488 -1577 -450
rect -1777 -505 -1727 -488
rect -1885 -522 -1869 -505
rect -2001 -538 -1869 -522
rect -1743 -522 -1727 -505
rect -1627 -505 -1577 -488
rect -1519 -488 -1319 -450
rect -1519 -505 -1469 -488
rect -1627 -522 -1611 -505
rect -1743 -538 -1611 -522
rect -1485 -522 -1469 -505
rect -1369 -505 -1319 -488
rect -1261 -488 -1061 -450
rect -1261 -505 -1211 -488
rect -1369 -522 -1353 -505
rect -1485 -538 -1353 -522
rect -1227 -522 -1211 -505
rect -1111 -505 -1061 -488
rect -1003 -488 -803 -450
rect -1003 -505 -953 -488
rect -1111 -522 -1095 -505
rect -1227 -538 -1095 -522
rect -969 -522 -953 -505
rect -853 -505 -803 -488
rect -745 -488 -545 -450
rect -745 -505 -695 -488
rect -853 -522 -837 -505
rect -969 -538 -837 -522
rect -711 -522 -695 -505
rect -595 -505 -545 -488
rect -487 -488 -287 -450
rect -487 -505 -437 -488
rect -595 -522 -579 -505
rect -711 -538 -579 -522
rect -453 -522 -437 -505
rect -337 -505 -287 -488
rect -229 -488 -29 -450
rect -229 -505 -179 -488
rect -337 -522 -321 -505
rect -453 -538 -321 -522
rect -195 -522 -179 -505
rect -79 -505 -29 -488
rect 29 -488 229 -450
rect 29 -505 79 -488
rect -79 -522 -63 -505
rect -195 -538 -63 -522
rect 63 -522 79 -505
rect 179 -505 229 -488
rect 287 -488 487 -450
rect 287 -505 337 -488
rect 179 -522 195 -505
rect 63 -538 195 -522
rect 321 -522 337 -505
rect 437 -505 487 -488
rect 545 -488 745 -450
rect 545 -505 595 -488
rect 437 -522 453 -505
rect 321 -538 453 -522
rect 579 -522 595 -505
rect 695 -505 745 -488
rect 803 -488 1003 -450
rect 803 -505 853 -488
rect 695 -522 711 -505
rect 579 -538 711 -522
rect 837 -522 853 -505
rect 953 -505 1003 -488
rect 1061 -488 1261 -450
rect 1061 -505 1111 -488
rect 953 -522 969 -505
rect 837 -538 969 -522
rect 1095 -522 1111 -505
rect 1211 -505 1261 -488
rect 1319 -488 1519 -450
rect 1319 -505 1369 -488
rect 1211 -522 1227 -505
rect 1095 -538 1227 -522
rect 1353 -522 1369 -505
rect 1469 -505 1519 -488
rect 1577 -488 1777 -450
rect 1577 -505 1627 -488
rect 1469 -522 1485 -505
rect 1353 -538 1485 -522
rect 1611 -522 1627 -505
rect 1727 -505 1777 -488
rect 1835 -488 2035 -450
rect 1835 -505 1885 -488
rect 1727 -522 1743 -505
rect 1611 -538 1743 -522
rect 1869 -522 1885 -505
rect 1985 -505 2035 -488
rect 2093 -488 2293 -450
rect 2093 -505 2143 -488
rect 1985 -522 2001 -505
rect 1869 -538 2001 -522
rect 2127 -522 2143 -505
rect 2243 -505 2293 -488
rect 2351 -488 2551 -450
rect 2351 -505 2401 -488
rect 2243 -522 2259 -505
rect 2127 -538 2259 -522
rect 2385 -522 2401 -505
rect 2501 -505 2551 -488
rect 2609 -488 2809 -450
rect 2609 -505 2659 -488
rect 2501 -522 2517 -505
rect 2385 -538 2517 -522
rect 2643 -522 2659 -505
rect 2759 -505 2809 -488
rect 2867 -488 3067 -450
rect 2867 -505 2917 -488
rect 2759 -522 2775 -505
rect 2643 -538 2775 -522
rect 2901 -522 2917 -505
rect 3017 -505 3067 -488
rect 3125 -488 3325 -450
rect 3125 -505 3175 -488
rect 3017 -522 3033 -505
rect 2901 -538 3033 -522
rect 3159 -522 3175 -505
rect 3275 -505 3325 -488
rect 3383 -488 3583 -450
rect 3383 -505 3433 -488
rect 3275 -522 3291 -505
rect 3159 -538 3291 -522
rect 3417 -522 3433 -505
rect 3533 -505 3583 -488
rect 3641 -488 3841 -450
rect 3641 -505 3691 -488
rect 3533 -522 3549 -505
rect 3417 -538 3549 -522
rect 3675 -522 3691 -505
rect 3791 -505 3841 -488
rect 3791 -522 3807 -505
rect 3675 -538 3807 -522
<< polycont >>
rect -3791 488 -3691 522
rect -3533 488 -3433 522
rect -3275 488 -3175 522
rect -3017 488 -2917 522
rect -2759 488 -2659 522
rect -2501 488 -2401 522
rect -2243 488 -2143 522
rect -1985 488 -1885 522
rect -1727 488 -1627 522
rect -1469 488 -1369 522
rect -1211 488 -1111 522
rect -953 488 -853 522
rect -695 488 -595 522
rect -437 488 -337 522
rect -179 488 -79 522
rect 79 488 179 522
rect 337 488 437 522
rect 595 488 695 522
rect 853 488 953 522
rect 1111 488 1211 522
rect 1369 488 1469 522
rect 1627 488 1727 522
rect 1885 488 1985 522
rect 2143 488 2243 522
rect 2401 488 2501 522
rect 2659 488 2759 522
rect 2917 488 3017 522
rect 3175 488 3275 522
rect 3433 488 3533 522
rect 3691 488 3791 522
rect -3791 -522 -3691 -488
rect -3533 -522 -3433 -488
rect -3275 -522 -3175 -488
rect -3017 -522 -2917 -488
rect -2759 -522 -2659 -488
rect -2501 -522 -2401 -488
rect -2243 -522 -2143 -488
rect -1985 -522 -1885 -488
rect -1727 -522 -1627 -488
rect -1469 -522 -1369 -488
rect -1211 -522 -1111 -488
rect -953 -522 -853 -488
rect -695 -522 -595 -488
rect -437 -522 -337 -488
rect -179 -522 -79 -488
rect 79 -522 179 -488
rect 337 -522 437 -488
rect 595 -522 695 -488
rect 853 -522 953 -488
rect 1111 -522 1211 -488
rect 1369 -522 1469 -488
rect 1627 -522 1727 -488
rect 1885 -522 1985 -488
rect 2143 -522 2243 -488
rect 2401 -522 2501 -488
rect 2659 -522 2759 -488
rect 2917 -522 3017 -488
rect 3175 -522 3275 -488
rect 3433 -522 3533 -488
rect 3691 -522 3791 -488
<< locali >>
rect -4021 626 -3925 660
rect 3925 626 4021 660
rect -4021 564 -3987 626
rect 3987 564 4021 626
rect -3807 488 -3791 522
rect -3691 488 -3675 522
rect -3549 488 -3533 522
rect -3433 488 -3417 522
rect -3291 488 -3275 522
rect -3175 488 -3159 522
rect -3033 488 -3017 522
rect -2917 488 -2901 522
rect -2775 488 -2759 522
rect -2659 488 -2643 522
rect -2517 488 -2501 522
rect -2401 488 -2385 522
rect -2259 488 -2243 522
rect -2143 488 -2127 522
rect -2001 488 -1985 522
rect -1885 488 -1869 522
rect -1743 488 -1727 522
rect -1627 488 -1611 522
rect -1485 488 -1469 522
rect -1369 488 -1353 522
rect -1227 488 -1211 522
rect -1111 488 -1095 522
rect -969 488 -953 522
rect -853 488 -837 522
rect -711 488 -695 522
rect -595 488 -579 522
rect -453 488 -437 522
rect -337 488 -321 522
rect -195 488 -179 522
rect -79 488 -63 522
rect 63 488 79 522
rect 179 488 195 522
rect 321 488 337 522
rect 437 488 453 522
rect 579 488 595 522
rect 695 488 711 522
rect 837 488 853 522
rect 953 488 969 522
rect 1095 488 1111 522
rect 1211 488 1227 522
rect 1353 488 1369 522
rect 1469 488 1485 522
rect 1611 488 1627 522
rect 1727 488 1743 522
rect 1869 488 1885 522
rect 1985 488 2001 522
rect 2127 488 2143 522
rect 2243 488 2259 522
rect 2385 488 2401 522
rect 2501 488 2517 522
rect 2643 488 2659 522
rect 2759 488 2775 522
rect 2901 488 2917 522
rect 3017 488 3033 522
rect 3159 488 3175 522
rect 3275 488 3291 522
rect 3417 488 3433 522
rect 3533 488 3549 522
rect 3675 488 3691 522
rect 3791 488 3807 522
rect -3887 438 -3853 454
rect -3887 -454 -3853 -438
rect -3629 438 -3595 454
rect -3629 -454 -3595 -438
rect -3371 438 -3337 454
rect -3371 -454 -3337 -438
rect -3113 438 -3079 454
rect -3113 -454 -3079 -438
rect -2855 438 -2821 454
rect -2855 -454 -2821 -438
rect -2597 438 -2563 454
rect -2597 -454 -2563 -438
rect -2339 438 -2305 454
rect -2339 -454 -2305 -438
rect -2081 438 -2047 454
rect -2081 -454 -2047 -438
rect -1823 438 -1789 454
rect -1823 -454 -1789 -438
rect -1565 438 -1531 454
rect -1565 -454 -1531 -438
rect -1307 438 -1273 454
rect -1307 -454 -1273 -438
rect -1049 438 -1015 454
rect -1049 -454 -1015 -438
rect -791 438 -757 454
rect -791 -454 -757 -438
rect -533 438 -499 454
rect -533 -454 -499 -438
rect -275 438 -241 454
rect -275 -454 -241 -438
rect -17 438 17 454
rect -17 -454 17 -438
rect 241 438 275 454
rect 241 -454 275 -438
rect 499 438 533 454
rect 499 -454 533 -438
rect 757 438 791 454
rect 757 -454 791 -438
rect 1015 438 1049 454
rect 1015 -454 1049 -438
rect 1273 438 1307 454
rect 1273 -454 1307 -438
rect 1531 438 1565 454
rect 1531 -454 1565 -438
rect 1789 438 1823 454
rect 1789 -454 1823 -438
rect 2047 438 2081 454
rect 2047 -454 2081 -438
rect 2305 438 2339 454
rect 2305 -454 2339 -438
rect 2563 438 2597 454
rect 2563 -454 2597 -438
rect 2821 438 2855 454
rect 2821 -454 2855 -438
rect 3079 438 3113 454
rect 3079 -454 3113 -438
rect 3337 438 3371 454
rect 3337 -454 3371 -438
rect 3595 438 3629 454
rect 3595 -454 3629 -438
rect 3853 438 3887 454
rect 3853 -454 3887 -438
rect -3807 -522 -3791 -488
rect -3691 -522 -3675 -488
rect -3549 -522 -3533 -488
rect -3433 -522 -3417 -488
rect -3291 -522 -3275 -488
rect -3175 -522 -3159 -488
rect -3033 -522 -3017 -488
rect -2917 -522 -2901 -488
rect -2775 -522 -2759 -488
rect -2659 -522 -2643 -488
rect -2517 -522 -2501 -488
rect -2401 -522 -2385 -488
rect -2259 -522 -2243 -488
rect -2143 -522 -2127 -488
rect -2001 -522 -1985 -488
rect -1885 -522 -1869 -488
rect -1743 -522 -1727 -488
rect -1627 -522 -1611 -488
rect -1485 -522 -1469 -488
rect -1369 -522 -1353 -488
rect -1227 -522 -1211 -488
rect -1111 -522 -1095 -488
rect -969 -522 -953 -488
rect -853 -522 -837 -488
rect -711 -522 -695 -488
rect -595 -522 -579 -488
rect -453 -522 -437 -488
rect -337 -522 -321 -488
rect -195 -522 -179 -488
rect -79 -522 -63 -488
rect 63 -522 79 -488
rect 179 -522 195 -488
rect 321 -522 337 -488
rect 437 -522 453 -488
rect 579 -522 595 -488
rect 695 -522 711 -488
rect 837 -522 853 -488
rect 953 -522 969 -488
rect 1095 -522 1111 -488
rect 1211 -522 1227 -488
rect 1353 -522 1369 -488
rect 1469 -522 1485 -488
rect 1611 -522 1627 -488
rect 1727 -522 1743 -488
rect 1869 -522 1885 -488
rect 1985 -522 2001 -488
rect 2127 -522 2143 -488
rect 2243 -522 2259 -488
rect 2385 -522 2401 -488
rect 2501 -522 2517 -488
rect 2643 -522 2659 -488
rect 2759 -522 2775 -488
rect 2901 -522 2917 -488
rect 3017 -522 3033 -488
rect 3159 -522 3175 -488
rect 3275 -522 3291 -488
rect 3417 -522 3433 -488
rect 3533 -522 3549 -488
rect 3675 -522 3691 -488
rect 3791 -522 3807 -488
rect -4021 -626 -3987 -564
rect 3987 -626 4021 -564
rect -4021 -660 -3925 -626
rect 3925 -660 4021 -626
<< viali >>
rect -3791 488 -3691 522
rect -3533 488 -3433 522
rect -3275 488 -3175 522
rect -3017 488 -2917 522
rect -2759 488 -2659 522
rect -2501 488 -2401 522
rect -2243 488 -2143 522
rect -1985 488 -1885 522
rect -1727 488 -1627 522
rect -1469 488 -1369 522
rect -1211 488 -1111 522
rect -953 488 -853 522
rect -695 488 -595 522
rect -437 488 -337 522
rect -179 488 -79 522
rect 79 488 179 522
rect 337 488 437 522
rect 595 488 695 522
rect 853 488 953 522
rect 1111 488 1211 522
rect 1369 488 1469 522
rect 1627 488 1727 522
rect 1885 488 1985 522
rect 2143 488 2243 522
rect 2401 488 2501 522
rect 2659 488 2759 522
rect 2917 488 3017 522
rect 3175 488 3275 522
rect 3433 488 3533 522
rect 3691 488 3791 522
rect -3887 -438 -3853 438
rect -3629 -438 -3595 438
rect -3371 -438 -3337 438
rect -3113 -438 -3079 438
rect -2855 -438 -2821 438
rect -2597 -438 -2563 438
rect -2339 -438 -2305 438
rect -2081 -438 -2047 438
rect -1823 -438 -1789 438
rect -1565 -438 -1531 438
rect -1307 -438 -1273 438
rect -1049 -438 -1015 438
rect -791 -438 -757 438
rect -533 -438 -499 438
rect -275 -438 -241 438
rect -17 -438 17 438
rect 241 -438 275 438
rect 499 -438 533 438
rect 757 -438 791 438
rect 1015 -438 1049 438
rect 1273 -438 1307 438
rect 1531 -438 1565 438
rect 1789 -438 1823 438
rect 2047 -438 2081 438
rect 2305 -438 2339 438
rect 2563 -438 2597 438
rect 2821 -438 2855 438
rect 3079 -438 3113 438
rect 3337 -438 3371 438
rect 3595 -438 3629 438
rect 3853 -438 3887 438
rect -3791 -522 -3691 -488
rect -3533 -522 -3433 -488
rect -3275 -522 -3175 -488
rect -3017 -522 -2917 -488
rect -2759 -522 -2659 -488
rect -2501 -522 -2401 -488
rect -2243 -522 -2143 -488
rect -1985 -522 -1885 -488
rect -1727 -522 -1627 -488
rect -1469 -522 -1369 -488
rect -1211 -522 -1111 -488
rect -953 -522 -853 -488
rect -695 -522 -595 -488
rect -437 -522 -337 -488
rect -179 -522 -79 -488
rect 79 -522 179 -488
rect 337 -522 437 -488
rect 595 -522 695 -488
rect 853 -522 953 -488
rect 1111 -522 1211 -488
rect 1369 -522 1469 -488
rect 1627 -522 1727 -488
rect 1885 -522 1985 -488
rect 2143 -522 2243 -488
rect 2401 -522 2501 -488
rect 2659 -522 2759 -488
rect 2917 -522 3017 -488
rect 3175 -522 3275 -488
rect 3433 -522 3533 -488
rect 3691 -522 3791 -488
<< metal1 >>
rect -3803 522 -3679 528
rect -3803 488 -3791 522
rect -3691 488 -3679 522
rect -3803 482 -3679 488
rect -3545 522 -3421 528
rect -3545 488 -3533 522
rect -3433 488 -3421 522
rect -3545 482 -3421 488
rect -3287 522 -3163 528
rect -3287 488 -3275 522
rect -3175 488 -3163 522
rect -3287 482 -3163 488
rect -3029 522 -2905 528
rect -3029 488 -3017 522
rect -2917 488 -2905 522
rect -3029 482 -2905 488
rect -2771 522 -2647 528
rect -2771 488 -2759 522
rect -2659 488 -2647 522
rect -2771 482 -2647 488
rect -2513 522 -2389 528
rect -2513 488 -2501 522
rect -2401 488 -2389 522
rect -2513 482 -2389 488
rect -2255 522 -2131 528
rect -2255 488 -2243 522
rect -2143 488 -2131 522
rect -2255 482 -2131 488
rect -1997 522 -1873 528
rect -1997 488 -1985 522
rect -1885 488 -1873 522
rect -1997 482 -1873 488
rect -1739 522 -1615 528
rect -1739 488 -1727 522
rect -1627 488 -1615 522
rect -1739 482 -1615 488
rect -1481 522 -1357 528
rect -1481 488 -1469 522
rect -1369 488 -1357 522
rect -1481 482 -1357 488
rect -1223 522 -1099 528
rect -1223 488 -1211 522
rect -1111 488 -1099 522
rect -1223 482 -1099 488
rect -965 522 -841 528
rect -965 488 -953 522
rect -853 488 -841 522
rect -965 482 -841 488
rect -707 522 -583 528
rect -707 488 -695 522
rect -595 488 -583 522
rect -707 482 -583 488
rect -449 522 -325 528
rect -449 488 -437 522
rect -337 488 -325 522
rect -449 482 -325 488
rect -191 522 -67 528
rect -191 488 -179 522
rect -79 488 -67 522
rect -191 482 -67 488
rect 67 522 191 528
rect 67 488 79 522
rect 179 488 191 522
rect 67 482 191 488
rect 325 522 449 528
rect 325 488 337 522
rect 437 488 449 522
rect 325 482 449 488
rect 583 522 707 528
rect 583 488 595 522
rect 695 488 707 522
rect 583 482 707 488
rect 841 522 965 528
rect 841 488 853 522
rect 953 488 965 522
rect 841 482 965 488
rect 1099 522 1223 528
rect 1099 488 1111 522
rect 1211 488 1223 522
rect 1099 482 1223 488
rect 1357 522 1481 528
rect 1357 488 1369 522
rect 1469 488 1481 522
rect 1357 482 1481 488
rect 1615 522 1739 528
rect 1615 488 1627 522
rect 1727 488 1739 522
rect 1615 482 1739 488
rect 1873 522 1997 528
rect 1873 488 1885 522
rect 1985 488 1997 522
rect 1873 482 1997 488
rect 2131 522 2255 528
rect 2131 488 2143 522
rect 2243 488 2255 522
rect 2131 482 2255 488
rect 2389 522 2513 528
rect 2389 488 2401 522
rect 2501 488 2513 522
rect 2389 482 2513 488
rect 2647 522 2771 528
rect 2647 488 2659 522
rect 2759 488 2771 522
rect 2647 482 2771 488
rect 2905 522 3029 528
rect 2905 488 2917 522
rect 3017 488 3029 522
rect 2905 482 3029 488
rect 3163 522 3287 528
rect 3163 488 3175 522
rect 3275 488 3287 522
rect 3163 482 3287 488
rect 3421 522 3545 528
rect 3421 488 3433 522
rect 3533 488 3545 522
rect 3421 482 3545 488
rect 3679 522 3803 528
rect 3679 488 3691 522
rect 3791 488 3803 522
rect 3679 482 3803 488
rect -3893 438 -3847 450
rect -3893 -438 -3887 438
rect -3853 -438 -3847 438
rect -3893 -450 -3847 -438
rect -3635 438 -3589 450
rect -3635 -438 -3629 438
rect -3595 -438 -3589 438
rect -3635 -450 -3589 -438
rect -3377 438 -3331 450
rect -3377 -438 -3371 438
rect -3337 -438 -3331 438
rect -3377 -450 -3331 -438
rect -3119 438 -3073 450
rect -3119 -438 -3113 438
rect -3079 -438 -3073 438
rect -3119 -450 -3073 -438
rect -2861 438 -2815 450
rect -2861 -438 -2855 438
rect -2821 -438 -2815 438
rect -2861 -450 -2815 -438
rect -2603 438 -2557 450
rect -2603 -438 -2597 438
rect -2563 -438 -2557 438
rect -2603 -450 -2557 -438
rect -2345 438 -2299 450
rect -2345 -438 -2339 438
rect -2305 -438 -2299 438
rect -2345 -450 -2299 -438
rect -2087 438 -2041 450
rect -2087 -438 -2081 438
rect -2047 -438 -2041 438
rect -2087 -450 -2041 -438
rect -1829 438 -1783 450
rect -1829 -438 -1823 438
rect -1789 -438 -1783 438
rect -1829 -450 -1783 -438
rect -1571 438 -1525 450
rect -1571 -438 -1565 438
rect -1531 -438 -1525 438
rect -1571 -450 -1525 -438
rect -1313 438 -1267 450
rect -1313 -438 -1307 438
rect -1273 -438 -1267 438
rect -1313 -450 -1267 -438
rect -1055 438 -1009 450
rect -1055 -438 -1049 438
rect -1015 -438 -1009 438
rect -1055 -450 -1009 -438
rect -797 438 -751 450
rect -797 -438 -791 438
rect -757 -438 -751 438
rect -797 -450 -751 -438
rect -539 438 -493 450
rect -539 -438 -533 438
rect -499 -438 -493 438
rect -539 -450 -493 -438
rect -281 438 -235 450
rect -281 -438 -275 438
rect -241 -438 -235 438
rect -281 -450 -235 -438
rect -23 438 23 450
rect -23 -438 -17 438
rect 17 -438 23 438
rect -23 -450 23 -438
rect 235 438 281 450
rect 235 -438 241 438
rect 275 -438 281 438
rect 235 -450 281 -438
rect 493 438 539 450
rect 493 -438 499 438
rect 533 -438 539 438
rect 493 -450 539 -438
rect 751 438 797 450
rect 751 -438 757 438
rect 791 -438 797 438
rect 751 -450 797 -438
rect 1009 438 1055 450
rect 1009 -438 1015 438
rect 1049 -438 1055 438
rect 1009 -450 1055 -438
rect 1267 438 1313 450
rect 1267 -438 1273 438
rect 1307 -438 1313 438
rect 1267 -450 1313 -438
rect 1525 438 1571 450
rect 1525 -438 1531 438
rect 1565 -438 1571 438
rect 1525 -450 1571 -438
rect 1783 438 1829 450
rect 1783 -438 1789 438
rect 1823 -438 1829 438
rect 1783 -450 1829 -438
rect 2041 438 2087 450
rect 2041 -438 2047 438
rect 2081 -438 2087 438
rect 2041 -450 2087 -438
rect 2299 438 2345 450
rect 2299 -438 2305 438
rect 2339 -438 2345 438
rect 2299 -450 2345 -438
rect 2557 438 2603 450
rect 2557 -438 2563 438
rect 2597 -438 2603 438
rect 2557 -450 2603 -438
rect 2815 438 2861 450
rect 2815 -438 2821 438
rect 2855 -438 2861 438
rect 2815 -450 2861 -438
rect 3073 438 3119 450
rect 3073 -438 3079 438
rect 3113 -438 3119 438
rect 3073 -450 3119 -438
rect 3331 438 3377 450
rect 3331 -438 3337 438
rect 3371 -438 3377 438
rect 3331 -450 3377 -438
rect 3589 438 3635 450
rect 3589 -438 3595 438
rect 3629 -438 3635 438
rect 3589 -450 3635 -438
rect 3847 438 3893 450
rect 3847 -438 3853 438
rect 3887 -438 3893 438
rect 3847 -450 3893 -438
rect -3803 -488 -3679 -482
rect -3803 -522 -3791 -488
rect -3691 -522 -3679 -488
rect -3803 -528 -3679 -522
rect -3545 -488 -3421 -482
rect -3545 -522 -3533 -488
rect -3433 -522 -3421 -488
rect -3545 -528 -3421 -522
rect -3287 -488 -3163 -482
rect -3287 -522 -3275 -488
rect -3175 -522 -3163 -488
rect -3287 -528 -3163 -522
rect -3029 -488 -2905 -482
rect -3029 -522 -3017 -488
rect -2917 -522 -2905 -488
rect -3029 -528 -2905 -522
rect -2771 -488 -2647 -482
rect -2771 -522 -2759 -488
rect -2659 -522 -2647 -488
rect -2771 -528 -2647 -522
rect -2513 -488 -2389 -482
rect -2513 -522 -2501 -488
rect -2401 -522 -2389 -488
rect -2513 -528 -2389 -522
rect -2255 -488 -2131 -482
rect -2255 -522 -2243 -488
rect -2143 -522 -2131 -488
rect -2255 -528 -2131 -522
rect -1997 -488 -1873 -482
rect -1997 -522 -1985 -488
rect -1885 -522 -1873 -488
rect -1997 -528 -1873 -522
rect -1739 -488 -1615 -482
rect -1739 -522 -1727 -488
rect -1627 -522 -1615 -488
rect -1739 -528 -1615 -522
rect -1481 -488 -1357 -482
rect -1481 -522 -1469 -488
rect -1369 -522 -1357 -488
rect -1481 -528 -1357 -522
rect -1223 -488 -1099 -482
rect -1223 -522 -1211 -488
rect -1111 -522 -1099 -488
rect -1223 -528 -1099 -522
rect -965 -488 -841 -482
rect -965 -522 -953 -488
rect -853 -522 -841 -488
rect -965 -528 -841 -522
rect -707 -488 -583 -482
rect -707 -522 -695 -488
rect -595 -522 -583 -488
rect -707 -528 -583 -522
rect -449 -488 -325 -482
rect -449 -522 -437 -488
rect -337 -522 -325 -488
rect -449 -528 -325 -522
rect -191 -488 -67 -482
rect -191 -522 -179 -488
rect -79 -522 -67 -488
rect -191 -528 -67 -522
rect 67 -488 191 -482
rect 67 -522 79 -488
rect 179 -522 191 -488
rect 67 -528 191 -522
rect 325 -488 449 -482
rect 325 -522 337 -488
rect 437 -522 449 -488
rect 325 -528 449 -522
rect 583 -488 707 -482
rect 583 -522 595 -488
rect 695 -522 707 -488
rect 583 -528 707 -522
rect 841 -488 965 -482
rect 841 -522 853 -488
rect 953 -522 965 -488
rect 841 -528 965 -522
rect 1099 -488 1223 -482
rect 1099 -522 1111 -488
rect 1211 -522 1223 -488
rect 1099 -528 1223 -522
rect 1357 -488 1481 -482
rect 1357 -522 1369 -488
rect 1469 -522 1481 -488
rect 1357 -528 1481 -522
rect 1615 -488 1739 -482
rect 1615 -522 1627 -488
rect 1727 -522 1739 -488
rect 1615 -528 1739 -522
rect 1873 -488 1997 -482
rect 1873 -522 1885 -488
rect 1985 -522 1997 -488
rect 1873 -528 1997 -522
rect 2131 -488 2255 -482
rect 2131 -522 2143 -488
rect 2243 -522 2255 -488
rect 2131 -528 2255 -522
rect 2389 -488 2513 -482
rect 2389 -522 2401 -488
rect 2501 -522 2513 -488
rect 2389 -528 2513 -522
rect 2647 -488 2771 -482
rect 2647 -522 2659 -488
rect 2759 -522 2771 -488
rect 2647 -528 2771 -522
rect 2905 -488 3029 -482
rect 2905 -522 2917 -488
rect 3017 -522 3029 -488
rect 2905 -528 3029 -522
rect 3163 -488 3287 -482
rect 3163 -522 3175 -488
rect 3275 -522 3287 -488
rect 3163 -528 3287 -522
rect 3421 -488 3545 -482
rect 3421 -522 3433 -488
rect 3533 -522 3545 -488
rect 3421 -528 3545 -522
rect 3679 -488 3803 -482
rect 3679 -522 3691 -488
rect 3791 -522 3803 -488
rect 3679 -528 3803 -522
<< properties >>
string FIXED_BBOX -4004 -643 4004 643
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.5 l 1 m 1 nf 30 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 60 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
